LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 1436; 
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00110" & "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000" & "111111111111111111000000000000000000011111111111110000000000000000000000000000011111111111111111000000000000000000001111111111111111000000011111111111111111000000000001111111111111111100000000000011111111111111111100000000000000000000001111111111111111110000000111111111111111111000000000000000111111111111111111000000000000000000000000111111111111111111000000011111111111111111100000000000000000000000111111111111111111000000000000000000111111111111000000000000000111111111111111110000000000000000011111111111111111100000000000000000000000000000111111111111111111000000000000000000111111111111111111000000000000000000000000001111111111111111100000000000000000000000000011111111111111111000000000000000011111111111111111100000000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000000000111111111111111111000000000000001111111111111111110000000001111111111111111110000000000000000001111111111111111100000000000000000000000001111111111111110000000000000000000000000000001111111111111111100000001111111111111111100000000000000000000000000000001111111111111110000000011111111111111111100000000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000111111111111111111000000000001111111111111111110000000000000000000000000000000111111111111111111000000000000000000000000000111111111111111111000000000000000000011111111111111111100000000000000000";
    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000" & "011001000100110110000000000000000000011111000110010000000000000000000000000000000101111101000011000000000000000000000010010111001011000000010101100011001001000000000001110110101110001000000000000000101100000110111100000000000000000000001010100001000110110000000111100111111100001000000000000000101011001110101001000000000000000000000000101001000011011000000000011100011010110100000000000000000000000000011000011111010100000000000000000000111000111011000000000000000011011000011010100000000000000000010101110100001010100000000000000000000000000000001101000101010100000000000000000000001010000100011111000000000000000000000000000010010010001000100000000000000000000000000010100101100011100000000000000000010111001101110111000000000000000000000000000000010000010100010100000000000000000000000010110110110001110000000000000000000000000000000001011000100001110000000000000001110011110010101000000000001110101111111110010000000000000000000011001001111001000000000000000000000000000010000111110100000000000000000000000000000000010110001010111000000001110011010111010100000000000000000000000000000001110000111100010000000010101010111010101000000000000000000000000000000010100001100111000000000000000000000000000010010000000011110000000000000000101101010001010001000000000001011111001101001000000000000000000000000000000000101011011010001110000000000000000000000000000001101000011110101000000000000000000000100100001110100100000000000000000";

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (  
				34 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				134 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				141 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				218 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				325 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				360 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				369 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				413 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				423 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				576 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				599 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				632 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				645 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				657 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				662 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				761 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				768 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				826 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				841 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				877 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				976 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				1105 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				1195 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				1225 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				1252 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				1281 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				1285 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				1359 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				1384 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				1433 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				1479 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				1490 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				1570 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				1586 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				1641 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				1666 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				1669 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				1784 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				1853 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				1934 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				1943 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				1946 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				2003 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				2051 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				2141 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				2153 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				2175 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				2182 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				2297 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				2444 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				2493 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				2497 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				2533 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				2585 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				2602 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				2670 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				2704 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				2732 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				2760 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				2867 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				2988 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				3040 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				3052 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				3066 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				3072 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				3087 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				3122 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				3156 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				3308 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				3311 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				3327 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				3328 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				3342 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				3377 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				3381 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				3429 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				3487 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				3495 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				3552 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				3595 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				3630 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				3667 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				3679 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				3700 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				3723 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				3730 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				3822 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				3827 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				3838 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				3849 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				3854 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				3868 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				3889 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				3904 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				3945 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				3986 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				4020 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				4021 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				4063 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				4081 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				4092 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				4116 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				4147 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				4167 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				4172 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				4231 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				4242 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				4265 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				4329 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				4371 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				4445 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				4501 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				4505 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				4519 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				4640 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				4667 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				4681 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				4697 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				4737 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				4756 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				4797 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				4806 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				4860 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				4888 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				4896 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				4908 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				4954 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				4984 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				5054 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				5056 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				5059 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				5062 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				5088 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				5089 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				5167 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				5198 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				5225 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				5288 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				5303 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				5329 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				5338 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				5348 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				5361 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				5363 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				5376 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				5390 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				5396 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				5487 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				5517 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				5573 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				5610 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				5614 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				5618 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				5624 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				5668 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				5869 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				5906 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				5954 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				6017 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				6085 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				6280 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				6307 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				6345 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				6353 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				6366 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				6379 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				6449 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				6473 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				6497 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				6523 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				6593 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				6701 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				6822 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				6902 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				6904 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				7092 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				7115 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				7137 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				7174 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				7179 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				7204 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				7236 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				7282 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				7285 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				7290 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				7314 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				7346 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				7369 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				7391 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				7488 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				7490 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				7520 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				7539 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				7586 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				7616 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				7652 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				7679 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				7680 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				7710 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				7731 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				7743 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				7748 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				7775 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				7811 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				7861 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				7880 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				8007 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				8014 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				8031 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				8056 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				8071 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				8091 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				8107 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				8160 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				8162 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				8179 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				8229 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				8240 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				8349 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				8364 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				8485 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				8496 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				8500 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				8533 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				8543 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				8563 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				8606 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				8640 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				8722 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				8725 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				8768 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				8839 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				8841 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				8860 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				8911 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				9015 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				9034 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				9035 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				9041 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				9054 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				9061 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				9083 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				9092 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				9099 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				9127 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				9184 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				9194 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				9196 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				9258 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				9279 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				9298 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				9333 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				9365 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				9409 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				9521 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				9568 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				9664 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				9666 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				9716 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				9757 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				9809 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				9830 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				9859 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				9921 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				9962 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				10008 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				10066 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				10070 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				10078 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				10085 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				10102 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				10159 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				10225 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				10226 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				10353 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				10356 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				10373 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				10384 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				10387 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				10461 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				10462 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				10467 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				10498 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				10523 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				10586 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				10615 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				10660 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				10730 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				10744 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				10798 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				10840 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				10852 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				10870 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				10893 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				10977 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				10988 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				11000 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				11079 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				11111 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				11151 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				11173 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				11190 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				11201 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				11226 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				11249 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				11315 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				11365 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				11403 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				11404 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				11468 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				11490 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				11501 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				11520 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				11600 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				11610 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				11675 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				11684 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				11769 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				11772 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				11916 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				11936 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				12015 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				12026 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				12091 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				12097 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				12153 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				12165 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				12168 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				12230 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				12266 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				12292 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				12300 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				12329 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				12352 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				12388 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				12412 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				12425 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				12426 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				12437 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				12459 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				12479 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				12499 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				12503 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				12528 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				12618 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				12644 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				12663 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				12671 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				12741 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				12798 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				12834 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				13005 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				13008 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				13028 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				13032 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				13078 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				13093 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				13099 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				13102 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				13191 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				13225 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				13277 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				13299 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				13316 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				13323 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				13351 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				13353 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				13388 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				13398 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				13460 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				13463 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				13479 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				13482 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				13550 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				13563 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				13630 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				13663 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				13666 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				13678 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				13692 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				13713 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				13759 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				13761 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				13768 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				13800 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				13879 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				13915 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				14024 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				14043 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				14068 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				14114 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				14124 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				14137 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				14138 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				14187 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				14233 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				14292 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				14356 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				14373 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				14394 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				14574 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				14577 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				14587 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				14702 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				14708 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				14734 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				14773 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				14831 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				14841 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				14872 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				14932 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				14952 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				14966 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				14969 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				14972 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				14974 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				14977 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				15006 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				15066 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				15074 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				15104 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				15150 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				15240 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				15317 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				15589 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				15602 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				15609 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				15614 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				15626 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				15645 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				15721 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				15730 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				15750 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				15757 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				15763 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				15911 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				16107 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				16148 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				16156 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				16158 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				16220 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				16256 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				16299 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				16352 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				16429 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				16443 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				16447 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				16491 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				16515 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				16604 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				16605 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				16639 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				16693 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				16704 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				16739 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				16765 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				16769 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				16790 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				16815 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				16855 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				16969 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				17095 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				17119 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				17141 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				17195 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				17215 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				17223 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				17259 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				17269 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				17288 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				17302 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				17320 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				17349 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				17394 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				17416 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				17491 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				17492 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				17534 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				17555 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				17575 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				17583 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				17646 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				17672 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				17849 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				17920 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				18009 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				18047 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				18068 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				18100 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				18120 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				18178 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				18214 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				18287 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				18292 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				18295 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				18305 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				18309 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				18332 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				18354 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				18444 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				18461 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				18513 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				18565 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				18636 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				18658 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				18703 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				18726 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				18756 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				18911 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				18974 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				19014 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				19050 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				19102 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				19180 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				19264 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				19327 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				19420 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				19431 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				19445 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				19485 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				19518 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				19579 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				19602 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				19612 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				19777 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				19805 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				19825 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				19830 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				19841 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				19909 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				19978 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				20006 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				20012 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				20112 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				20118 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				20153 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				20169 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				20206 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				20238 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				20261 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				20358 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				20360 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				20387 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				20439 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				20442 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				20456 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				20462 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				20474 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				20489 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				20499 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				20560 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				20562 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				20571 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				20616 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				20696 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				20699 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				20708 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				20749 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				20782 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				20819 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				20996 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				21014 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				21058 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				21075 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				21121 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				21127 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				21212 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				21218 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				21309 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				21424 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				21468 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				21470 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				21477 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				21485 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				21515 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				21544 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				21567 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				21592 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				21601 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				21607 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				21612 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				21636 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				21654 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				21657 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				21684 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				21690 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				21722 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				21735 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				21798 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				21800 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				21828 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				21832 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				21855 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				21863 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				21935 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				21937 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				21953 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				21987 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				21990 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				22041 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				22129 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				22176 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				22186 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				22256 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				22261 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				22272 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				22419 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				22454 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				22515 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				22521 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				22590 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				22616 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				22624 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				22641 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				22691 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				22806 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				22814 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				22902 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				22922 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				22936 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				22940 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				22979 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				22995 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				23043 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				23048 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				23066 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				23074 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				23131 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				23140 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				23143 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				23146 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				23153 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				23165 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				23200 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				23222 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				23279 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				23293 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				23333 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				23352 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				23410 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				23412 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				23438 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				23461 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				23494 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				23580 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				23617 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				23674 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				23689 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				23705 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				23781 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				23790 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				23793 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				23805 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				23912 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				23935 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				23936 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				23947 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				24030 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				24133 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				24175 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				24258 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				24337 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				24418 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				24439 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				24475 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				24541 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				24552 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				24576 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				24600 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				24685 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				24702 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				24791 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				24834 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				24862 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				24865 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				24872 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				24906 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				25056 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				25065 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				25109 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				25113 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				25121 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				25141 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				25217 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				25219 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				25251 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				25278 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				25283 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				25333 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				25343 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				25355 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				25356 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				25407 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				25468 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				25507 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				25522 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				25664 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				25686 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				25739 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				25766 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				25826 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				25827 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				25923 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				25945 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				25966 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				25987 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				25998 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				26040 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				26060 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				26064 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				26223 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				26244 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				26249 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				26288 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				26321 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				26350 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				26398 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				26405 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				26461 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				26485 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				26489 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				26490 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				26559 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				26583 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				26651 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				26691 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				26698 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				26715 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				26717 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				26721 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				26743 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				26746 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				26789 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				26827 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				26837 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				26853 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				26880 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				26915 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				26958 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				26974 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				26976 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				27025 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				27032 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				27138 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				27178 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				27193 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				27255 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				27270 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				27275 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				27331 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				27376 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				27379 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				27406 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				27423 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				27558 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				27567 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				27583 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				27614 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				27627 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				27672 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				27696 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				27725 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				27792 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				27804 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				27810 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				27879 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				27930 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				27942 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				27951 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				28081 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				28169 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				28207 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				28246 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				28256 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				28312 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				28356 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				28359 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				28366 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				28408 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				28415 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				28458 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				28535 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				28547 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				28589 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				28609 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				28618 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				28666 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				28688 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				28718 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				28727 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				28731 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				28737 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				28745 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				28833 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				28879 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				28934 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				28944 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				28997 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				28999 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				29006 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				29020 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				29085 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				29106 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				29177 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				29179 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				29204 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				29233 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				29235 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				29269 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				29304 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				29326 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				29358 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				29409 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				29446 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				29454 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				29460 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				29465 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				29531 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				29553 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				29655 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				29810 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				29914 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				29966 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				30016 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				30028 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				30110 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				30145 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				30160 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				30218 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				30258 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				30271 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				30291 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				30314 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				30362 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				30381 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				30460 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				30495 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				30501 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				30537 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				30541 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				30588 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				30595 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				30638 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				30652 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				30681 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				30731 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				30749 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				30756 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				30905 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				30953 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				30972 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				31023 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				31030 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				31038 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				31039 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				31056 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				31109 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				31228 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				31288 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				31300 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				31353 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				31431 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				31460 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				31541 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				31588 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				31624 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				31627 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				31688 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				31704 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				31799 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				31814 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				31841 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				31863 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				31891 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				31936 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				31956 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				31973 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				32111 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				32154 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				32235 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				32257 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				32282 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				32283 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				32321 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				32329 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				32413 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				32422 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				32449 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				32456 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				32474 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				32477 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				32514 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				32550 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				32662 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				32688 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				32692 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				32725 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				32733 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				32772 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				32821 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				32832 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				32996 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				33032 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				33049 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				33097 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				33103 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				33133 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				33152 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				33183 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				33189 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				33195 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				33198 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				33209 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				33242 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				33260 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				33261 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				33271 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				33328 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				33333 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				33351 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				33356 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				33374 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				33393 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				33404 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				33418 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				33445 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				33473 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				33513 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				33538 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				33548 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				33583 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				33618 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				33673 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				33681 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				33692 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				33748 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				33755 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				33772 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				33774 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				33855 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				33886 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				33936 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				33949 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				33981 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				34020 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				34043 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				34081 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				34090 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				34103 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				34177 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				34211 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				34235 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				34241 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				34256 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				34316 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				34336 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				34474 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				34591 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				34620 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				34639 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				34669 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				34672 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				34673 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				34690 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				34715 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				34748 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				34782 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				34798 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				34812 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				34874 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				34900 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				34931 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				34977 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				35027 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				35060 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				35101 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				35136 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				35194 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				35245 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				35310 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				35337 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				35356 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				35369 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				35377 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				35393 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				35464 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				35467 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				35470 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				35478 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				35532 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				35561 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				35618 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				35644 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				35651 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				35722 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				35815 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				35838 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				35862 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				35865 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				35907 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				35926 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				36055 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				36063 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				36123 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				36145 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				36152 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				36176 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				36235 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				36284 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				36294 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				36335 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				36358 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				36363 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				36372 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				36408 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				36441 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				36465 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				36502 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				36594 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				36600 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				36626 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				36722 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				36760 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				36796 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				36797 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				36800 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				36803 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				36816 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				36870 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				36880 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				36972 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				36976 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				36989 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				37075 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				37081 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				37138 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				37141 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				37186 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				37205 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				37293 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				37341 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				37367 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				37377 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				37409 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				37414 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				37569 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				37591 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				37596 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				37660 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				37690 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				37748 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				37765 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				37800 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				37845 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				37895 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				37920 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				37960 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				38021 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				38044 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				38122 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				38148 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				38169 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				38272 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				38297 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				38299 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				38358 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				38361 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				38367 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				38403 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				38454 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				38585 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				38626 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				38632 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				38676 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				38759 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				38862 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				38870 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				38881 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				38937 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				38950 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				38960 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				39042 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				39057 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				39060 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				39076 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				39212 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				39255 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				39265 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				39276 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				39284 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				39317 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				39387 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				39432 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				39449 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				39476 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				39500 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				39520 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				39570 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				39605 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				39615 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				39644 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				39668 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				39736 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				39750 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				39753 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				39756 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				39771 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				39810 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				39841 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				39976 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				40026 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				40036 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				40069 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				40132 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				40196 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				40248 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				40256 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				40284 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				40299 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				40337 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				40355 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				40439 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				40443 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				40466 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				40504 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				40521 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				40577 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				40617 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				40623 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				40683 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				40717 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				40724 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				40750 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				40849 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				40869 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				40873 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				40896 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				40925 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				40930 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				40971 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				41015 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				41048 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				41062 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				41080 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				41188 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				41201 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				41287 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				41306 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				41311 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				41312 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				41346 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				41371 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				41377 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				41383 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				41438 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				41458 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				41496 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				41509 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				41578 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				41591 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				41698 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				41737 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				41738 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				41752 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				41810 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				41825 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				41827 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				41880 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				41895 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				41900 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				41935 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				41954 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				42025 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				42038 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				42048 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				42109 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				42122 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				42199 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				42229 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				42239 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				42310 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				42335 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				42394 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				42406 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				42458 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				42474 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				42528 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				42547 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				42554 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				42624 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				42632 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				42685 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				42712 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				42757 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				42860 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				43001 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				43029 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				43040 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				43049 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				43196 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				43214 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				43261 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				43275 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				43281 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				43318 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				43365 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				43397 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				43401 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				43469 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				43519 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				43556 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				43564 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				43598 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				43671 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				43691 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				43728 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				43742 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				43766 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				43774 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				43777 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				43838 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				43887 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				43899 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				43911 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				43944 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				44009 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				44034 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				44047 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				44063 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				44080 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				44082 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				44125 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				44126 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				44137 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				44142 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				44198 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				44210 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				44212 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				44228 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				44257 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				44325 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				44355 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				44408 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				44409 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				44426 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				44441 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				44472 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				44575 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				44662 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				44671 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				44691 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				44723 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				44838 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				44854 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				44887 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				44901 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				44948 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				44982 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				45021 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				45050 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				45067 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				45103 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				45121 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				45154 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				45155 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				45175 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				45233 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				45236 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				45249 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				45518 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				45524 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				45587 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				45627 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				45702 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				45757 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				45778 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				45807 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				45818 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				45846 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				45875 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				45943 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				46000 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				46062 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				46068 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				46079 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				46085 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				46171 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				46227 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				46322 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				46387 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				46411 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				46422 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				46451 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				46485 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				46558 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				46591 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				46594 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				46604 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				46618 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				46631 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				46671 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				46697 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				46839 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				46857 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				46872 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				46928 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				46975 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				47004 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				47006 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				47068 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				47107 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				47129 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				47163 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				47185 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				47230 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				47277 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				47286 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				47290 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				47347 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				47357 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				47363 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				47440 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				47443 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				47495 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				47508 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				47545 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				47617 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				47688 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				47757 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				47778 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				47784 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				47819 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				47895 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				47912 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				47918 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				47924 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				47938 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				48097 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				48111 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				48145 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				48175 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				48237 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				48288 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				48292 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				48308 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				48320 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				48325 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				48355 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				48413 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				48437 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				48472 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				48478 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				48513 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				48516 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				48580 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				48599 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				48715 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				48720 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				48822 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				48864 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				48890 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				48982 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				49013 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				49024 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				49040 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				49067 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				49080 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				49096 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				49109 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				49295 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				49353 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				49388 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				49408 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				49477 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				49572 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				49703 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				49716 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				49739 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				49757 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				49779 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				49822 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				49826 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				49879 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				49915 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				49930 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				49974 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				50033 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				50089 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				50090 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				50207 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				50265 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				50283 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				50288 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				50308 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				50311 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				50317 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				50328 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				50330 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				50331 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				50346 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				50424 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				50491 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				50523 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				50532 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				50587 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				50651 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				50695 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				50743 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				50746 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				50753 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				50878 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				50981 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				51017 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				51095 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				51137 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				51152 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				51159 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				51169 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				51222 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				51279 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				51288 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				51314 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				51395 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				51431 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				51439 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				51461 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				51517 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				51523 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				51537 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				51540 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				51543 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				51627 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				51649 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				51673 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				51691 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				51748 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				51817 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				51853 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				51856 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				51918 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				51923 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				51926 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				52013 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				52043 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				52069 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				52112 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				52138 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				52195 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				52207 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				52238 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				52244 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				52266 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				52270 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				52317 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				52343 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				52392 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				52396 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				52408 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				52429 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				52446 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				52518 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				52528 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				52693 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				52727 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				52743 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				52747 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				52773 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				52775 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				52788 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				52805 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				52862 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				52885 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				52968 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				52977 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				52990 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				52996 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				52999 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				53009 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				53020 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				53091 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				53116 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				53130 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				53134 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				53193 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				53212 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				53240 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				53285 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				53337 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				53340 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				53413 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				53456 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				53484 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				53562 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				53618 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				53622 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				53626 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				53628 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				53634 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				53661 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				53726 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				53749 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				53779 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				53792 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				53840 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				53849 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				53901 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				53979 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				54052 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				54078 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				54096 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				54097 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				54132 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				54177 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				54193 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				54243 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				54265 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				54305 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				54317 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				54379 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				54382 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				54386 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				54402 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				54454 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				54456 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				54605 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				54611 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				54672 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				54782 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				54789 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				54814 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				54841 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				54843 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				54853 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				54861 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				54876 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				54888 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				54895 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				54919 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				54954 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				54972 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				54983 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				55000 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				55007 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				55061 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				55140 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				55264 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				55432 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				55449 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				55487 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				55508 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				55538 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				55596 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				55633 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				55641 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				55647 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				55649 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				55659 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				55661 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				55662 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				55671 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				55695 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				55702 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				55750 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				55798 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				55963 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				55968 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				55978 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				56027 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				56126 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				56127 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				56157 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				56170 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				56233 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				56291 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				56430 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				56463 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				56506 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				56511 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				56555 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				56606 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				56625 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				56673 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				56745 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				56751 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				56788 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				56816 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				56882 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				56887 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				56964 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				57017 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				57036 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				57087 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				57132 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				57133 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				57153 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				57200 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				57210 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				57244 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				57275 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				57308 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				57313 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				57316 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				57334 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				57342 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				57405 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				57417 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				57477 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				57575 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				57579 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				57598 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				57617 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				57665 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				57728 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				57779 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				57849 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				57878 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				57912 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				57940 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				57953 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				57977 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				57995 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				58049 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				58083 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				58109 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				58117 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				58129 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				58144 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				58196 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				58203 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				58223 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				58245 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				58250 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				58272 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				58290 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				58315 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				58331 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				58369 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				58389 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				58517 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				58546 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				58570 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				58574 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				58587 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				58634 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				58657 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				58670 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				58731 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				58786 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				58789 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				58793 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				58813 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				58846 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				58958 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				58978 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				59000 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				59010 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				59031 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				59112 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				59121 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				59131 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				59154 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				59183 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				59188 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				59194 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				59213 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				59239 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				59419 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				59460 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				59468 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				59474 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				59549 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				59554 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				59603 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				59639 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				59658 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				59681 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				59715 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				59731 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				59738 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				59779 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				59933 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				60009 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				60061 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				60221 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				60302 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				60338 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				60361 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				60413 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				60428 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				60452 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				60525 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				60527 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				60531 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				60559 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				60635 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				60642 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				60664 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				60717 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				60733 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				60807 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				60836 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				60861 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				60935 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				61083 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				61143 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				61152 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				61176 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				61243 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				61245 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				61258 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				61302 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				61404 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				61436 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				61519 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				61567 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				61653 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				61654 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				61680 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				61772 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				61781 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				61852 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				61869 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				62055 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				62062 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				62089 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				62096 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				62167 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				62319 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				62412 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				62437 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				62463 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				62530 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				62542 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				62566 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				62571 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				62590 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				62604 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				62638 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				62662 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				62700 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				62757 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				62786 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				62788 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				62811 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				62823 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				62848 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				62929 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				62932 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				62980 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				62987 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				63013 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				63024 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				63040 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				63110 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				63174 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				63217 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				63258 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				63275 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				63320 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				63380 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				63396 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				63397 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				63448 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				63466 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				63542 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				63582 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				63599 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				63606 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				63638 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				63667 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				63747 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				63760 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				63928 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				63930 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				63981 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				64038 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				64050 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				64074 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				64188 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				64200 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				64211 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				64229 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				64280 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				64294 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				64451 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				64470 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				64478 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				64566 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				64567 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				64575 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				64692 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				64714 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				64770 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				64871 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				64896 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				64934 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				64946 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				65009 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				65123 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				65136 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				65161 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				65162 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				65233 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				65272 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				65284 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				65334 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				65392 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				65419 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				65476 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),

                                OTHERS => STD_LOGIC_VECTOR(to_unsigned(240, 8))
                            );
                    
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
                ASSERT (mem_we = '1' OR mem_we = '0') REPORT "o_mem_we in an unexpected state" SEVERITY failure;
            END IF;
            ASSERT (enable_wire = '1' OR enable_wire = '0') REPORT "o_mem_en in an unexpected state" SEVERITY failure;
        END IF;
    END PROCESS;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    createScenario : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '0' THEN
            tb_rst <= scenario_rst(0);
            tb_w <= scenario_w(0);
            tb_start <= scenario_start(0);
            scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_done = '0' REPORT "TEST FALLITO (postreset DONE != 0 )" SEVERITY failure;
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1001000100110110:240->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 11100011001:240->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 101111101000011:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 10010111001011:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 101100011001001:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 101101011100010:240->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1011000001101111:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1010000100011011:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1100111111100001:240->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1011001110101001:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1001000011011000:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1000110101101000:240->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1000011111010100:240->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1000111011:240->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 101100001101010:240->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1011101000010101:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1101000101010100:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1010000100011111:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 100100100010001:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 100101100011100:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1110011011101110:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(154, 8)) severity failure; -- 1000001010001010:154->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(154, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1101101100011100:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1011000100001110:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1001111001010100:240->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1010111111111001:240->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 110010011110010:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1000011111010:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 101100010101110:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 100110101110101:240->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1000011110001:240->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1010101110101010:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 100001100111000:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1001000000001111:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1101010001010001:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1111100110100100:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1011011010001110:240->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1101000011110101:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- 1001000011101001:240->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 

        ASSERT false REPORT "Simulation Ended! TEST PASSATO (EXAMPLE)" SEVERITY failure;
    END PROCESS testRoutine;

END projecttb;