LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 2748; 
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00110" & "0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000" & "1111111111111111110000000000000000000000000001111111111111111110000000000001111111111111111110000000000011111111111111111000000000000000111111111111111111000111111111111111111000000000000000000001111111111111111110000000000000000000011111111111100000000000000000001111111111111111000000000000000000000000001111111111111000001111111111111111100000000000000000000000000000011111111111111111100000000000000011111111111111000000000000000000011111111111111111100000000000000000000000000000111111111111000011111111111111111100000000000000000000000000011111111111110000000000000000000011111111111111110000000000000001111111111111111110000000011111111111111111000000000000000000000000000011111111111111111101111111111111111000000000000000000111111111111111110000000000000000000000000011111111111111111100000000000000000000000000000111111111111111111000000000111111111111111111000011111111111111110000000000000000000000000000001111111111111111000000000000000000000000000000111111111111111111000000000000000000011111111111111110000000000000111111111111111110000000000000000000001111111111111111110000111111111111111110000000000000000000000000001111111111111111110000000000000000000000000000000111111111111111111000000000000000000000000001111111111111111100000000000000000011111111111111111100000000000000000000000011111111111111111000000000001111111111111111110000000000000000000011111111111111111001111111111111111100000000000000000000000000001111111111111111100000000000000000000001111111111111111100001111111111111111100000000011111111111111111000000000000000000000000111111111111111111000000111111111111111111000000000000000000000000001111111111111000000000000000011111111111111111000000000000000001111111111111111110000000000000000000000000000011111111111111111000000000000011111111000000000000000000000000011111111111111111000000000011111111111111111100000000000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000011111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000111111111111111111000000000001111111111111000000000000000000000000000000011111111111111111100011111111111111100000000111111111111110000000000000111111111111111000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111110000000000000000111111111111111111000000000000000000000000111111111111111100000111111111111111110000000000000000001111111111111111000000000000000000000000000111111111111111111000000000000000000111111111111111111000000000000000000000000000111111111111111100000000000000000000000000000111111111111100000000000000000001111111111111111100000111111111111111111000000000000001111111111111111110011111111111111100000000000000000000000";
    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000" & "1100110101100010110000000000000000000000000000111010001011101010000000000001100101000101100010000000000011111010001111011000000000000000011000110001111001000011111011000011111000000000000000000000101010110101000110000000000000000000011100111111100000000000000000001011011000111111000000000000000000000000001011000100001000001000011100111110100000000000000000000000000000010111000010111100100000000000000011111000001101000000000000000000000111110000011101100000000000000000000000000000000111011111000000101011110100010100000000000000000000000000001011110001110000000000000000000000110110011010010000000000000000110011110001100010000000000101110011011001000000000000000000000000000011010000100110111100001111010111111000000000000000000001010110011110110000000000000000000000000010010011110011001100000000000000000000000000000101010010010001101000000000001001100011110001000010101010001001010000000000000000000000000000000111010011011011000000000000000000000000000000101000000100011001000000000000000000000100110101010010000000000000001001001001101010000000000000000000000010000111000000010000101101111110011010000000000000000000000000000001011010011101110000000000000000000000000000000010101001100110101000000000000000000000000001100101101100000100000000000000000001100101101100001100000000000000000000000010001011110011111000000000000000110110100100110000000000000000000010101100100011111000101011110001000100000000000000000000000000001110110110111100100000000000000000000000011101110000011100001001110110101111100000000011001100110011011000000000000000000000000110100101110101001000000010101011010001101000000000000000000000000000100001001001000000000000000000000000101010001000000000000000000100110111010011010000000000000000000000000000011110001010000011000000000000001100101000000000000000000000000001101110110010101000000000001001111010000100100000000000000000000000000000001011111111111011010000000000000000000000000001001010100101110100000010110100100010000000000000000000000000011000111100000101000000000000000000000111100011000001111000000000000010010101001100011000000000001011000001101000000000000000000000000000000010001000001000111100011001001100110100000000101111101101110000000000000100110101111001000000001000100111000001110000000000000000000000011100000000100110000000000000000000000001111010001110110000000000000000110000111011011101000000000000000000000000000010011010001100000110100111001101110000000000000000001001100001111001000000000000000000000000000101011100010100101000000000000000000110111101001010111000000000000000000000000000110111111011000100000000000000000000000000000000000110000100000000000000000001100101000110001100000100101101000000111000000000000001011001110110100110010010011000000100000000000000000000000";

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (  
				1 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				42 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				123 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				164 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				257 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				349 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				428 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				479 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				511 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				625 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				627 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				696 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				829 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				836 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				885 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				983 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				1166 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				1223 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				1304 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				1460 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				1510 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				1591 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				1613 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				1631 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				1652 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				1661 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				1759 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				1769 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				1853 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				1878 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				1902 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				1916 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				1937 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				1990 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				2064 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				2067 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				2208 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				2220 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				2230 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				2236 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				2238 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				2319 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				2420 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				2426 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				2477 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				2636 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				2649 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				2739 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				2839 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				3023 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				3071 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				3079 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				3162 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				3350 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				3376 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				3425 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				3432 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				3484 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				3495 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				3539 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				3642 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				3719 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				3758 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				3828 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				3850 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				4117 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				4124 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				4251 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				4257 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				4303 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				4376 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				4547 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				4579 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				4586 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				4608 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				4716 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				4739 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				4779 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				4783 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				4844 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				4853 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				4857 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				4910 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				5001 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				5031 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				5064 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				5094 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				5188 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				5190 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				5198 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				5272 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				5406 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				5415 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				5490 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				5499 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				5577 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				5698 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				5714 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				5796 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				5798 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				6060 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				6084 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				6227 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				6309 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				6330 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				6345 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				6456 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				6494 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				6497 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				6592 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				6593 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				6629 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				6703 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				6822 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				6842 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				6857 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				6910 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				6993 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				7034 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				7053 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				7072 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				7119 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				7134 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				7142 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				7147 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				7183 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				7222 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				7364 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				7396 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				7400 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				7407 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				7425 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				7479 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				7487 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				7548 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				7579 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				7689 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				7695 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				7753 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				7779 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				7789 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				7868 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				7877 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				7888 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				7909 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				7927 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				8012 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				8044 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				8195 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				8206 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				8225 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				8336 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				8464 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				8475 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				8528 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				8580 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				8782 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				8913 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				8950 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				8956 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				9032 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				9042 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				9046 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				9089 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				9133 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				9285 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				9296 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				9354 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				9375 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				9386 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				9426 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				9587 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				9693 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				9726 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				9790 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				9791 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				9871 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				10071 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				10138 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				10190 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				10213 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				10312 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				10360 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				10457 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				10605 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				10648 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				10695 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				10705 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				10727 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				10852 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				10889 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				10933 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				11048 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				11218 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				11338 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				11518 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				11544 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				11609 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				11677 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				11736 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				11737 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				11777 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				11967 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				11973 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				12018 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				12027 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				12038 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				12192 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				12226 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				12280 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				12316 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				12395 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				12429 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				12435 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				12491 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				12517 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				12540 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				12580 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				12614 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				12630 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				12676 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				12729 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				12815 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				12852 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				12865 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				12935 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				13017 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				13065 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				13133 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				13145 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				13204 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				13243 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				13309 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				13382 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				13419 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				13446 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				13454 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				13462 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				13532 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				13556 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				13581 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				13759 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				13788 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				13813 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				13828 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				13959 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				13968 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				14023 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				14048 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				14084 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				14130 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				14151 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				14189 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				14255 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				14325 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				14398 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				14408 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				14511 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				14631 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				14648 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				14700 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				14719 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				14736 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				14880 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				14925 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				14936 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				14938 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				14952 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				14988 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				15033 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				15111 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				15144 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				15145 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				15148 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				15198 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				15286 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				15329 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				15478 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				15494 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				15594 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				15621 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				15625 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				15707 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				15749 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				15752 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				15918 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				15928 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				15938 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				16017 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				16032 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				16117 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				16133 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				16287 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				16310 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				16324 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				16357 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				16437 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				16454 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				16609 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				16614 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				16626 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				16655 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				16657 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				16712 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				16767 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				16972 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				17064 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				17080 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				17083 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				17201 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				17215 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				17228 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				17380 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				17472 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				17537 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				17579 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				17586 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				17604 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				17650 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				17658 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				17659 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				17705 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				17897 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				17899 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				17908 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				17986 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				17988 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				17996 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				18003 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				18012 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				18016 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				18163 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				18167 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				18314 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				18335 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				18402 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				18456 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				18653 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				18655 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				18733 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				18761 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				18775 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				18945 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				19152 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				19195 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				19206 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				19292 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				19403 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				19425 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				19458 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				19496 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				19540 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				19579 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				19594 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				19631 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				19680 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				19721 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				19790 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				19798 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				19846 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				19896 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				20015 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				20046 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				20054 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				20110 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				20120 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				20125 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				20130 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				20159 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				20200 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				20208 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				20259 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				20312 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				20411 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				20452 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				20453 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				20484 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				20486 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				20579 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				20641 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				20660 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				20710 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				20776 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				20799 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				20808 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				20811 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				20823 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				20885 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				20950 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				21008 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				21217 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				21227 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				21319 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				21347 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				21351 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				21437 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				21463 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				21499 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				21551 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				21589 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				21622 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				21661 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				21775 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				21971 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				22020 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				22059 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				22195 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				22279 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				22323 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				22336 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				22462 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				22529 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				22569 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				22784 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				22835 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				22901 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				22910 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				23026 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				23064 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				23098 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				23152 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				23174 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				23222 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				23331 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				23367 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				23495 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				23654 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				23665 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				23706 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				23718 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				23730 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				23752 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				23776 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				23812 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				23846 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				23885 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				23903 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				23905 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				23917 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				23961 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				24020 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				24227 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				24320 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				24323 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				24336 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				24357 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				24360 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				24367 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				24461 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				24480 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				24547 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				24548 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				24558 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				24566 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				24688 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				24746 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				24768 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				24773 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				24819 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				24828 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				24850 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				25021 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				25044 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				25066 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				25138 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				25238 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				25259 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				25308 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				25381 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				25499 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				25597 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				25608 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				25700 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				25780 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				25840 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				25869 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				25914 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				26052 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				26081 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				26233 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				26256 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				26438 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				26462 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				26526 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				26641 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				26716 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				26738 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				26746 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				26773 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				26788 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				26864 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				26976 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				27075 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				27161 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				27217 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				27287 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				27320 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				27339 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				27389 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				27429 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				27436 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				27451 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				27543 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				27596 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				27616 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				27651 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				27683 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				27747 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				27752 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				27895 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				27922 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				28019 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				28030 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				28089 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				28155 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				28175 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				28228 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				28232 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				28256 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				28301 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				28336 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				28424 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				28447 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				28471 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				28542 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				28545 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				28622 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				28745 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				28835 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				28957 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				28993 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				29110 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				29156 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				29163 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				29197 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				29203 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				29233 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				29239 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				29286 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				29368 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				29471 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				29512 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				29552 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				29592 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				29615 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				29629 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				29666 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				29708 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				29714 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				29841 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				29884 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				30091 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				30143 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				30228 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				30345 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				30482 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				30524 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				30538 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				30541 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				30560 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				30605 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				30752 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				30855 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				30882 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				30916 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				30942 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				30976 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				31186 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				31567 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				31587 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				31597 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				31648 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				31718 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				31818 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				31966 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				32000 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				32038 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				32128 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				32177 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				32185 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				32186 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				32229 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				32315 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				32324 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				32368 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				32391 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				32409 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				32413 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				32456 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				32473 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				32498 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				32538 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				32563 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				32761 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				32788 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				32801 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				32829 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				32909 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				32987 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				33116 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				33136 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				33170 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				33334 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				33359 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				33365 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				33371 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				33419 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				33715 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				33803 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				33842 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				34201 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				34250 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				34268 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				34332 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				34350 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				34435 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				34558 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				34638 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				34666 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				34673 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				34682 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				34704 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				34756 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				34814 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				34836 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				34923 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				35009 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				35048 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				35119 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				35129 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				35149 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				35187 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				35284 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				35300 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				35344 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				35449 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				35520 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				35533 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				35598 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				35602 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				35696 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				35757 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				35758 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				35786 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				35914 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				35927 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				36012 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				36053 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				36057 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				36084 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				36256 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				36294 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				36299 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				36371 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				36376 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				36404 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				36411 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				36424 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				36442 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				36451 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				36542 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				36628 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				36642 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				36705 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				36712 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				36723 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				36725 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				36779 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				36815 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				36965 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				37003 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				37010 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				37048 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				37134 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				37175 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				37248 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				37304 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				37352 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				37447 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				37501 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				37536 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				37538 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				37566 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				37672 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				37699 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				37727 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				37746 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				37840 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				37863 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				37868 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				37876 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				37979 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				37991 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				37999 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				38019 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				38028 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				38045 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				38049 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				38097 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				38221 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				38224 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				38259 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				38292 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				38366 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				38390 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				38519 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				38543 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				38571 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				38639 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				38775 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				38777 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				38867 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				38876 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				38887 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				38965 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				38984 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				39100 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				39134 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				39245 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				39247 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				39286 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				39332 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				39336 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				39344 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				39557 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				39586 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				39602 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				39839 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				39858 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				39867 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				39965 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				40073 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				40088 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				40146 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				40172 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				40225 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				40264 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				40330 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				40336 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				40349 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				40359 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				40567 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				40758 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				40828 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				40832 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				40836 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				40940 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				40953 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				40958 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				40981 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				41034 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				41076 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				41083 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				41234 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				41243 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				41268 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				41269 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				41465 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				41632 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				41788 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				41908 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				41990 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				42062 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				42063 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				42099 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				42229 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				42260 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				42265 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				42267 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				42296 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				42346 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				42374 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				42381 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				42420 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				42451 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				42505 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				42599 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				42669 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				42758 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				42761 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				42794 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				42814 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				42860 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				43007 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				43176 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				43216 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				43270 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				43279 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				43361 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				43677 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				43769 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				43770 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				43842 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				43872 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				43901 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				43972 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				44144 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				44200 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				44303 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				44380 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				44402 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				44413 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				44457 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				44537 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				44568 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				44616 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				44708 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				44754 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				44761 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				44762 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				44861 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				44867 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				44879 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				44933 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				44937 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				44956 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				45009 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				45051 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				45112 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				45156 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				45203 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				45207 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				45275 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				45396 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				45419 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				45511 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				45542 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				45552 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				45573 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				45623 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				45851 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				45925 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				46022 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				46055 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				46082 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				46147 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				46314 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				46321 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				46348 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				46451 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				46456 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				46498 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				46546 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				46652 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				46703 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				46802 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				46830 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				46912 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				46940 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				47039 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				47115 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				47140 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				47142 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				47222 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				47343 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				47371 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				47403 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				47413 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				47484 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				47505 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				47562 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				47572 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				47574 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				47602 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				47711 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				47750 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				47783 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				47868 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				47929 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				47957 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				48008 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				48014 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				48149 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				48173 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				48312 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				48339 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				48342 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				48452 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				48527 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				48596 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				48624 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				48641 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				48646 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				48711 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				48828 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				48882 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				48919 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				48940 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				48993 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				49066 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				49087 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				49125 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				49244 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				49365 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				49373 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				49506 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				49518 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				49573 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				49587 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				49654 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				49662 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				49801 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				49872 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				49919 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				49983 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				50036 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				50101 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				50132 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				50159 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				50168 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				50189 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				50191 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				50294 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				50323 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				50327 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				50359 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				50404 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				50451 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				50539 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				50659 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				50675 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				50792 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				50803 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				50833 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				50851 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				50859 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				50909 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				50967 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				50975 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				51035 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				51101 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				51152 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				51312 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				51318 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				51326 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				51458 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				51527 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				51539 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				51582 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				51598 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				51616 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				51641 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				51654 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				51657 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				51711 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				51786 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				51861 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				51865 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				51927 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				51948 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				52036 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				52048 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				52108 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				52259 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				52281 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				52304 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				52323 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				52346 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				52393 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				52416 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				52542 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				52559 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				52580 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				52649 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				52651 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				52886 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				52914 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				52935 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				52958 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				52960 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				53146 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				53159 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				53307 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				53416 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				53417 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				53476 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				53569 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				53628 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				53632 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				53660 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				53691 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				53908 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				53930 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				53959 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				54042 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				54111 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				54114 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				54145 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				54151 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				54176 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				54265 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				54388 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				54489 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				54646 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				54772 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				54906 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				54908 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				54962 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				55041 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				55096 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				55104 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				55123 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				55135 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				55219 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				55221 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				55239 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				55257 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				55277 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				55297 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				55363 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				55370 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				55372 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				55435 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				55450 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				55473 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				55525 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				55531 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				55613 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				55661 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				55711 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				55729 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				55740 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				55761 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				55777 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				55814 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				55878 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				55907 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				55917 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				55975 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				55987 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				56030 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				56127 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				56162 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				56172 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				56179 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				56314 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				56343 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				56687 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				56706 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				56770 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				56807 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				56812 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				56903 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				57013 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				57140 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				57146 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				57149 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				57197 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				57269 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				57286 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				57402 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				57406 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				57422 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				57450 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				57459 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				57469 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				57537 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				57592 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				57651 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				57673 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				57674 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				57900 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				57932 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				57954 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				58010 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				58015 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				58071 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				58163 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				58378 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				58398 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				58416 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				58445 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				58495 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				58588 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				58734 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				58888 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				58889 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				58894 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				58916 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				58955 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				58972 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				59021 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				59042 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				59147 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				59149 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				59182 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				59298 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				59511 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				59774 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				59872 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				59890 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				59919 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				59949 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				60012 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				60081 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				60089 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				60133 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				60148 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				60194 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				60274 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				60334 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				60421 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				60470 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				60591 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				60617 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				60654 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				60700 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				60832 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				60885 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				60912 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				60924 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				60984 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				61031 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				61076 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				61121 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				61249 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				61265 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				61277 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				61290 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				61320 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				61403 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				61415 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				61499 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				61540 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				61547 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				61552 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				61600 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				61777 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				61779 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				61818 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				61840 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				62038 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				62105 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				62160 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				62178 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				62179 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				62212 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				62233 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				62287 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				62297 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				62389 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				62460 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				62538 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				62553 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				62768 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				62770 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				62782 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				62864 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				62921 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				63018 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				63024 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				63187 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				63241 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				63242 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				63256 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				63266 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				63295 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				63304 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				63330 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				63365 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				63605 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				63693 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				63710 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				63982 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				64098 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				64108 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				64193 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				64231 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				64313 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				64432 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				64472 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				64551 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				64571 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				64622 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				64713 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				64734 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				64766 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				64788 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				64809 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				64824 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				64837 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				64864 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				65054 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				65060 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				65083 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				65153 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				65267 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				65313 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				65360 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				65413 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				65482 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				65500 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),

                                OTHERS => STD_LOGIC_VECTOR(to_unsigned(11, 8)
                            );
                    
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
                ASSERT (mem_we = '1' OR mem_we = '0') REPORT "o_mem_we in an unexpected state" SEVERITY failure;
            END IF;
            ASSERT (enable_wire = '1' OR enable_wire = '0') REPORT "o_mem_en in an unexpected state" SEVERITY failure;
        END IF;
    END PROCESS;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    createScenario : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '0' THEN
            tb_rst <= scenario_rst(0);
            tb_w <= scenario_w(0);
            tb_start <= scenario_start(0);
            scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_done = '0' REPORT "TEST FALLITO (postreset DONE != 0 )" SEVERITY failure;
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0011010110001011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1101000101110101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0010100010110001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --111010001111011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1000110001111001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1111011000011111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0101011010100011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1001111111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --11011000111111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --11000100001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --000111001111101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1110000101111001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --111000001101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1111100000111011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0111011111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1010111101000101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --01111000111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --11011001101001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1001111000110001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --101110011011001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0100001001101111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --01111010111111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --101011001111011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0100111100110011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1010010010001101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1001100011110001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --10101000100101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --11010011011011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1000000100011001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --10011010101001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --100100100110101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1000011100000001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --110111111001101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0101101001110111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0101001100110101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --001011011000001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1001011011000011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --001011110011111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0011011010010011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --101100100011111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --010111100010001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --101101101111001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --111011100000111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --011101101011111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --001100110011011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0100101110101001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0101011010001101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --00001001001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --000000101010001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0011011101001101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --110001010000011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --100101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --101110110010101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0011110100001001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1111111111101101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0010101001011101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --11010010001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1000111100000101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1100011000001111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0010101001100011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --11000001101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0010000010001111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0010011001101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --111110110111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0110101111001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0010011100000111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(11, 8)) severity failure; --110000000010011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1101000111011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0000111011011101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --00100110100011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --010011100110111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --01100001111001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1011100010100101:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0111101001010111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --01111110110001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8)) severity failure; --00001100001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8)) severity failure; --001010001100011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0101101000000111:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --1100111011010011:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8)) severity failure; --0100110000001:11
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 

        ASSERT false REPORT "Simulation Ended! TEST PASSATO (EXAMPLE)" SEVERITY failure;
    END PROCESS testRoutine;

END projecttb;