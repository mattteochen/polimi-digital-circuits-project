LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 1369; 
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00110" & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000" & "11111111111111000000000000000000000000111111111111111110000000000000000000000000001111111111111111110000000000000001111111111111111110000000000111111111111111111111111111111111110000000000000000111111111111111000000001111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111100000001111111111111111110000011111111000000000000000000011111111111100000000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000111111111111111000000000000001111111111111110000000001111111111111111100000000000000000000000000011111111111111110000000000000000001111111111111111100000000000000000111111111111111110000000000000000111111111111111111000000000000000000000001111111111111110000000011111111111111111100001111111111111111100000000000000001111111111111111100011111111111111111100000000000000000111111111111111111000000000000011111111111111111100000011111111111111110000001111111111111111110000000000000011111111111111111100001111111111111111100000000000000111111111111111110011111111111111111000000000000000000000000111111111111111111001111111111111111110000000000000000000000000000001111111111111111110000000000000111111111111111100000000000000000";
    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000" & "11110001011011000000000000000000000000111101011110001010000000000000000000000000001111110011011011110000000000000001101101001011000010000000000010110010000011110111000111100001110000000000000000011100111111111000000000010000100110110000000000000000000000000110110100110111100000000000000000000010101110111100101000000000000000000000000111110011000110100000001111011010010001110000001000001000000000000000000001001101110100000000000000000000000000000100110100100111000000000000000000000001111010110010110100000000000000000000001010110000011100010000000000000000000000001001010010100100000000000000000000010010011110001110100000000000000000101101001101111000000000000001010000010110010000000001001101111011011100000000000000000000000000001010100010100010000000000000000001001000110000100100000000000000000010100001000000110000000000000000101110011101010101000000000000000000000000100010110011110000000001100100011101001100000000010000010010100000000000000001011111111001100100011001100110001011100000000000000000011010001010111111000000000000010110111111111101100000010111101111101010000001000000000011101010000000000000000000110010110100100000001101011011101100000000000000011110000110101110011100101010110001000000000000000000000000011110111011111111000000101011011110010000000000000000000000000000000100010011011110110000000000000110001110111110100000000000000000";

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (  
				19 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				23 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				85 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				100 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				101 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				102 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				122 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				124 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				186 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				212 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				250 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				342 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				404 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				421 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				451 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				482 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				528 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				564 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				594 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				644 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				661 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				678 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				754 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				775 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				787 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				797 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				811 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				824 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				838 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				839 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				841 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				889 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				913 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				945 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				1071 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				1107 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				1129 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				1131 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				1133 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				1149 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				1172 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				1192 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				1206 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				1213 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				1272 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				1287 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				1343 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				1388 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				1422 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				1436 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				1480 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				1599 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				1612 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				1619 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				1631 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				1644 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				1745 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				1750 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				1765 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				1789 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				1819 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				1823 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				1862 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				1914 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				1917 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				1938 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				1945 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				2027 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				2059 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				2083 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				2110 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				2113 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				2125 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				2213 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				2277 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				2381 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				2383 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				2387 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				2398 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				2452 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				2467 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				2542 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				2596 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				2597 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				2598 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				2616 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				2628 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				2736 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				2790 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				2807 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				2862 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				2929 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				3042 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				3063 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				3086 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				3128 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				3150 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				3227 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				3300 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				3345 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				3433 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				3474 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				3511 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				3513 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				3557 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				3592 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				3632 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				3653 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				3740 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				3760 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				3768 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				3782 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				3799 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				3833 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				3840 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				3887 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				3889 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				3890 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				3909 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				3919 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				3921 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				3929 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				4078 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				4112 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				4165 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				4170 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				4206 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				4217 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				4239 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				4273 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				4335 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				4356 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				4380 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				4414 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				4437 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				4524 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				4526 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				4572 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				4579 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				4649 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				4664 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				4683 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				4752 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				4801 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				4836 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				4915 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				4919 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				4965 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				4971 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				5025 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				5030 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				5094 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				5144 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				5169 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				5171 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				5219 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				5281 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				5286 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				5299 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				5346 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				5352 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				5385 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				5387 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				5390 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				5484 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				5492 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				5506 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				5557 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				5594 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				5606 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				5687 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				5712 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				5805 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				5865 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				5886 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				5921 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				5999 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				6085 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				6165 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				6232 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				6319 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				6424 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				6426 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				6462 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				6481 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				6503 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				6516 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				6523 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				6530 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				6602 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				6635 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				6648 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				6686 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				6750 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				6768 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				6828 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				6841 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				6881 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				6904 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				6923 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				6928 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				6929 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				7020 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				7031 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				7085 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				7096 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				7130 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				7170 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				7237 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				7276 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				7291 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				7322 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				7424 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				7464 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				7485 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				7524 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				7577 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				7661 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				7662 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				7698 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				7709 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				7714 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				7757 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				7775 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				7787 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				7833 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				7841 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				7843 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				7877 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				7959 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				7961 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				8123 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				8210 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				8262 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				8276 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				8288 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				8300 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				8412 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				8416 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				8449 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				8468 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				8476 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				8495 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				8625 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				8638 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				8644 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				8722 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				8727 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				8729 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				8751 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				8753 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				8774 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				8942 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				9012 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				9022 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				9104 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				9143 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				9189 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				9229 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				9246 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				9252 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				9280 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				9324 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				9343 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				9353 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				9370 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				9388 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				9409 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				9437 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				9525 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				9528 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				9529 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				9604 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				9610 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				9626 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				9686 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				9839 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				9897 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				9908 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				9924 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				9974 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				10002 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				10023 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				10042 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				10049 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				10080 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				10143 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				10213 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				10226 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				10231 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				10236 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				10248 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				10258 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				10313 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				10332 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				10389 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				10393 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				10456 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				10485 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				10489 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				10497 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				10523 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				10561 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				10569 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				10643 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				10724 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				10756 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				10759 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				10817 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				10865 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				10866 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				10903 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				10971 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				10998 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				11000 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				11062 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				11095 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				11127 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				11195 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				11197 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				11267 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				11293 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				11301 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				11304 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				11325 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				11329 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				11385 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				11406 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				11474 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				11530 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				11599 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				11609 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				11612 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				11613 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				11627 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				11639 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				11768 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				11834 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				11850 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				11852 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				11950 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				12057 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				12104 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				12162 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				12179 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				12234 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				12296 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				12327 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				12338 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				12339 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				12439 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				12491 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				12726 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				12734 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				12774 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				12810 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				12890 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				12929 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				12939 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				12948 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				12950 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				12998 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				13003 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				13025 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				13067 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				13172 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				13184 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				13186 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				13204 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				13229 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				13265 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				13280 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				13282 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				13287 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				13351 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				13356 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				13372 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				13383 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				13400 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				13420 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				13430 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				13474 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				13477 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				13494 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				13518 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				13609 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				13629 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				13649 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				13674 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				13888 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				13893 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				13947 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				13985 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				13992 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				14029 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				14036 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				14126 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				14131 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				14132 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				14157 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				14186 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				14208 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				14241 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				14311 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				14324 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				14376 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				14421 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				14441 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				14468 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				14477 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				14493 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				14497 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				14519 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				14546 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				14614 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				14628 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				14638 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				14646 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				14730 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				14733 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				14820 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				14888 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				14910 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				14942 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				15011 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				15018 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				15025 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				15027 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				15048 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				15071 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				15103 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				15154 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				15178 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				15218 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				15227 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				15253 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				15285 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				15372 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				15401 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				15409 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				15431 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				15477 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				15520 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				15546 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				15550 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				15560 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				15570 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				15599 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				15669 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				15736 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				15757 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				15765 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				15769 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				15777 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				15780 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				15812 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				15834 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				15884 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				15891 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				15897 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				15902 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				15911 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				15961 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				16001 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				16031 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				16076 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				16093 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				16135 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				16170 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				16182 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				16187 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				16215 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				16256 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				16431 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				16451 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				16452 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				16455 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				16518 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				16632 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				16762 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				16793 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				16813 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				16829 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				16835 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				16877 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				16888 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				16971 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				16976 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				17035 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				17099 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				17131 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				17169 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				17237 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				17249 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				17260 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				17266 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				17289 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				17326 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				17347 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				17381 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				17389 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				17400 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				17441 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				17467 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				17497 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				17528 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				17540 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				17543 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				17573 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				17580 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				17600 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				17652 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				17662 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				17671 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				17689 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				17692 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				17719 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				17747 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				17762 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				17793 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				17857 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				17867 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				17914 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				17985 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				18016 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				18029 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				18039 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				18062 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				18131 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				18168 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				18170 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				18192 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				18207 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				18267 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				18307 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				18366 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				18409 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				18546 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				18555 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				18669 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				18675 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				18699 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				18755 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				18780 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				18883 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				18905 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				18923 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				19066 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				19147 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				19326 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				19330 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				19371 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				19375 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				19383 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				19442 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				19469 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				19478 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				19583 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				19602 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				19729 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				19743 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				19839 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				19846 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				19891 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				19961 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				20017 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				20065 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				20198 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				20230 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				20231 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				20278 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				20347 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				20348 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				20383 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				20389 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				20434 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				20451 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				20461 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				20542 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				20557 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				20569 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				20570 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				20590 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				20632 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				20639 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				20660 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				20713 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				20787 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				20816 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				20854 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				20908 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				20928 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				20974 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				20978 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				20985 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				21015 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				21021 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				21103 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				21188 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				21198 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				21215 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				21237 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				21282 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				21296 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				21297 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				21302 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				21303 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				21337 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				21401 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				21450 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				21510 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				21519 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				21546 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				21576 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				21626 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				21721 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				21726 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				21778 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				21806 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				21851 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				21862 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				21879 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				21939 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				21953 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				21973 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				21975 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				22047 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				22115 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				22136 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				22183 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				22214 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				22215 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				22269 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				22315 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				22396 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				22398 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				22412 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				22677 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				22686 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				22749 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				22751 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				22754 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				22768 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				22856 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				22866 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				22920 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				22982 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				23030 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				23063 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				23087 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				23102 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				23115 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				23300 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				23377 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				23388 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				23451 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				23475 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				23526 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				23536 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				23543 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				23613 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				23621 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				23643 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				23689 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				23692 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				23708 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				23734 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				23776 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				23816 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				23847 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				23968 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				24006 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				24033 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				24034 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				24155 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				24174 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				24192 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				24293 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				24296 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				24329 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				24331 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				24342 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				24433 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				24454 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				24493 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				24500 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				24503 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				24561 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				24581 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				24651 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				24666 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				24697 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				24698 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				24734 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				24747 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				24752 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				24775 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				24802 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				24880 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				24903 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				24988 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				25020 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				25042 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				25065 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				25317 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				25343 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				25387 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				25408 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				25414 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				25448 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				25460 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				25463 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				25493 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				25513 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				25522 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				25616 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				25696 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				25704 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				25727 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				25737 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				25837 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				25848 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				25856 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				25897 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				25943 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				26002 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				26067 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				26083 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				26112 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				26172 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				26197 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				26286 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				26432 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				26464 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				26495 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				26551 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				26569 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				26656 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				26660 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				26682 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				26719 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				26751 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				26986 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				27011 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				27018 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				27022 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				27036 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				27051 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				27091 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				27136 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				27262 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				27308 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				27467 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				27469 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				27533 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				27574 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				27584 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				27629 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				27753 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				27899 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				27934 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				28011 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				28064 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				28080 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				28168 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				28191 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				28248 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				28258 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				28394 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				28404 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				28420 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				28540 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				28567 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				28601 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				28642 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				28769 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				28800 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				28833 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				28835 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				28901 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				29043 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				29082 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				29105 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				29153 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				29177 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				29182 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				29223 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				29308 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				29326 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				29339 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				29382 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				29385 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				29419 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				29488 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				29511 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				29521 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				29630 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				29650 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				29698 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				29702 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				29779 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				29800 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				29844 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				29852 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				29899 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				29996 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				30017 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				30036 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				30058 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				30071 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				30135 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				30166 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				30219 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				30256 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				30257 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				30277 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				30304 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				30361 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				30423 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				30472 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				30532 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				30549 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				30631 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				30663 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				30682 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				30686 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				30692 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				30709 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				30765 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				30772 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				30777 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				30781 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				30794 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				30824 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				30885 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				30933 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				30971 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				30985 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				31057 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				31166 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				31173 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				31295 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				31303 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				31337 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				31347 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				31413 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				31493 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				31559 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				31580 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				31582 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				31612 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				31621 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				31672 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				31691 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				31724 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				31748 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				31759 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				31787 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				31826 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				31865 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				31884 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				31919 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				31949 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				31955 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				32026 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				32126 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				32138 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				32156 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				32162 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				32173 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				32182 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				32191 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				32202 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				32265 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				32316 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				32344 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				32442 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				32447 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				32460 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				32471 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				32499 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				32608 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				32610 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				32616 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				32631 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				32660 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				32688 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				32746 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				32758 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				32768 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				32786 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				32826 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				32854 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				32934 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				32997 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				33003 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				33144 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				33173 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				33217 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				33372 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				33384 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				33403 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				33448 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				33525 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				33529 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				33533 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				33536 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				33560 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				33615 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				33646 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				33676 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				33715 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				33800 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				33802 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				33890 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				33983 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				34019 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				34074 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				34185 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				34216 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				34247 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				34284 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				34380 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				34408 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				34437 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				34458 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				34556 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				34557 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				34587 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				34642 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				34767 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				34780 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				34786 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				34807 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				34808 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				34841 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				34879 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				34903 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				35049 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				35069 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				35080 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				35099 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				35202 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				35209 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				35255 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				35303 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				35331 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				35473 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				35551 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				35650 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				35663 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				35667 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				35724 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				35730 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				35735 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				35737 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				35748 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				35759 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				35796 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				35859 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				35871 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				35902 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				35936 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				36067 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				36109 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				36114 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				36138 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				36165 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				36198 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				36221 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				36245 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				36270 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				36319 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				36402 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				36405 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				36418 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				36503 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				36626 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				36630 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				36715 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				36754 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				36766 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				36793 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				36831 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				36860 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				36864 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				36865 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				36886 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				36907 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				36931 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				36986 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				36991 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				37025 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				37029 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				37046 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				37062 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				37090 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				37115 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				37180 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				37211 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				37215 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				37317 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				37338 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				37403 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				37442 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				37463 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				37541 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				37546 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				37599 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				37727 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				37746 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				37761 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				37787 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				37789 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				37800 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				37846 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				37888 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				37963 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				38027 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				38067 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				38119 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				38189 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				38220 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				38353 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				38367 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				38374 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				38381 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				38383 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				38432 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				38550 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				38681 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				38707 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				38715 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				38805 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				38816 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				38850 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				38954 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				38969 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				39076 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				39203 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				39204 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				39211 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				39218 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				39291 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				39329 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				39330 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				39331 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				39374 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				39456 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				39462 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				39471 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				39483 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				39557 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				39592 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				39596 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				39639 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				39673 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				39676 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				39712 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				39734 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				39911 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				39998 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				40063 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				40065 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				40079 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				40159 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				40163 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				40167 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				40169 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				40205 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				40221 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				40223 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				40274 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				40292 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				40312 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				40355 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				40407 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				40442 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				40523 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				40526 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				40645 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				40651 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				40667 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				40689 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				40695 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				40762 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				40769 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				40774 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				40827 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				40828 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				40844 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				40878 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				40884 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				40886 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				40940 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				40947 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				40952 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				40958 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				40971 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				40992 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				41019 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				41076 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				41176 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				41199 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				41242 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				41243 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				41247 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				41324 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				41344 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				41372 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				41550 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				41565 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				41572 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				41634 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				41745 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				41752 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				41772 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				41828 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				41936 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				41948 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				41970 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				41976 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				42019 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				42109 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				42137 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				42245 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				42273 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				42287 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				42321 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				42372 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				42373 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				42379 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				42394 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				42526 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				42566 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				42583 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				42587 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				42613 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				42632 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				42637 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				42641 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				42649 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				42739 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				42835 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				42849 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				42856 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				42901 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				42907 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				42951 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				42964 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				42971 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				43008 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				43048 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				43060 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				43088 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				43107 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				43122 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				43124 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				43150 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				43153 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				43218 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				43240 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				43255 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				43284 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				43334 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				43346 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				43356 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				43388 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				43472 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				43482 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				43518 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				43541 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				43561 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				43640 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				43654 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				43666 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				43671 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				43694 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				43699 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				43721 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				43742 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				43755 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				43795 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				43953 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				44026 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				44105 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				44117 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				44142 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				44151 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				44198 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				44258 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				44374 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				44406 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				44451 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				44497 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				44534 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				44535 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				44540 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				44593 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				44631 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				44650 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				44751 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				44825 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				44921 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				44974 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				44998 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				45083 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				45084 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				45109 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				45156 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				45193 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				45316 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				45322 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				45334 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				45384 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				45417 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				45431 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				45485 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				45488 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				45595 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				45597 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				45598 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				45611 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				45645 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				45661 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				45663 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				45682 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				45699 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				45713 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				45748 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				45758 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				45792 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				45911 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				45925 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				45937 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				45941 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				45952 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				45979 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				45985 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				46019 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				46060 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				46108 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				46136 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				46142 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				46155 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				46189 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				46196 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				46309 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				46311 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				46368 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				46385 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				46443 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				46491 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				46498 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				46520 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				46558 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				46584 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				46586 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				46634 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				46699 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				46702 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				46735 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				46811 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				46898 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				46938 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				47000 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				47018 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				47036 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				47042 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				47044 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				47092 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				47115 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				47117 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				47219 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				47318 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				47324 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				47395 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				47433 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				47453 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				47527 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				47536 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				47550 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				47555 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				47557 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				47569 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				47658 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				47676 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				47746 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				47763 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				47769 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				47783 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				47907 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				47931 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				47974 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				48089 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				48130 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				48190 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				48285 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				48291 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				48314 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				48401 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				48434 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				48482 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				48522 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				48535 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				48588 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				48603 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				48664 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				48665 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				48702 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				48766 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				48779 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				48780 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				48804 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				48807 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				48832 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				48855 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				48884 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				49051 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				49059 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				49154 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				49285 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				49293 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				49317 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				49324 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				49381 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				49391 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				49501 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				49560 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				49612 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				49627 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				49649 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				49730 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				49738 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				49750 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				49759 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				49823 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				49851 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				49856 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				49882 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				49894 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				49900 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				49907 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				49931 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				49985 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				50003 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				50035 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				50083 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				50098 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				50114 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				50120 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				50137 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				50145 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				50157 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				50169 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				50203 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				50210 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				50256 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				50272 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				50327 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				50349 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				50380 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				50411 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				50417 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				50427 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				50482 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				50544 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				50631 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				50773 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				50826 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				50843 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				50845 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				50893 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				50895 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				50911 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				50943 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				50967 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				51048 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				51071 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				51079 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				51163 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				51184 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				51196 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				51203 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				51246 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				51349 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				51352 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				51412 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				51420 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				51436 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				51524 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				51547 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				51559 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				51583 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				51704 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				51728 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				51756 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				51823 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				51831 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				51859 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				51985 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				51988 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				51992 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				52011 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				52092 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				52109 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				52162 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				52164 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				52174 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				52224 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				52237 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				52276 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				52297 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				52328 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				52382 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				52398 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				52399 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				52441 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				52469 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				52479 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				52490 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				52493 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				52499 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				52506 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				52512 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				52540 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				52603 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				52609 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				52705 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				52772 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				52788 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				52822 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				52834 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				52846 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				52848 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				52967 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				52993 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				53003 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				53058 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				53148 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				53225 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				53241 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				53298 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				53386 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				53404 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				53424 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				53429 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				53446 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				53468 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				53474 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				53479 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				53570 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				53603 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				53607 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				53631 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				53643 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				53646 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				53674 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				53725 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				53808 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				53824 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				53885 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				53922 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				53951 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				53961 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				54013 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				54051 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				54073 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				54121 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				54143 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				54154 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				54162 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				54188 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				54292 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				54312 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				54369 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				54456 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				54472 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				54499 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				54513 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				54514 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				54531 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				54576 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				54612 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				54730 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				54741 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				54771 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				54820 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				54838 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				54851 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				54855 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				54932 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				55005 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				55092 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				55095 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				55107 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				55113 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				55156 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				55230 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				55261 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				55275 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				55279 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				55297 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				55347 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				55355 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				55441 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				55549 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				55606 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				55613 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				55767 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				55769 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				55781 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				55951 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				55990 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				56135 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				56136 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				56149 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				56289 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				56294 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				56327 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				56366 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				56373 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				56401 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				56467 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				56516 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				56554 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				56566 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				56579 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				56598 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				56632 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				56731 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				56741 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				56759 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				56770 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				56798 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				56809 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				56834 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				56851 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				56883 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				56897 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				56988 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				57025 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				57042 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				57057 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				57078 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				57087 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				57093 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				57098 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				57152 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				57166 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				57186 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				57194 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				57258 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				57260 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				57261 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				57263 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				57301 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				57307 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				57331 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				57337 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				57348 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				57377 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				57388 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				57411 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				57537 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				57661 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				57668 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				57736 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				57856 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				57866 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				57983 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				58070 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				58092 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				58102 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				58115 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				58141 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				58185 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				58229 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				58246 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				58273 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				58295 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				58382 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				58399 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				58426 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				58441 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				58596 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				58705 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				58756 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				58807 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				58889 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				58930 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				58981 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				59004 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				59021 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				59116 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				59140 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				59184 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				59342 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				59392 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				59411 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				59469 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				59585 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				59625 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				59643 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				59663 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				59818 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				60009 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				60102 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				60151 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				60172 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				60189 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				60226 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				60265 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				60274 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				60346 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				60387 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				60428 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				60442 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				60490 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				60510 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				60520 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				60525 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				60559 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				60566 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				60623 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				60654 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				60656 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				60676 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				60737 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				60751 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				60769 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				60781 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				60792 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				60834 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				60858 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				60925 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				60933 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				60990 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				61003 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				61025 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				61052 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				61094 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				61107 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				61167 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				61192 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				61202 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				61221 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				61344 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				61401 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				61403 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				61442 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				61526 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				61588 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				61603 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				61660 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				61678 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				61688 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				61691 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				61834 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				61859 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				61894 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				61896 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				61919 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				61996 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				62034 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				62047 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				62079 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				62102 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				62139 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				62145 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				62295 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				62354 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				62456 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				62605 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				62635 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				62648 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				62652 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				62706 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				62751 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				62897 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				62923 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				62984 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				63028 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				63060 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				63099 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				63119 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				63122 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				63136 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				63158 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				63160 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				63259 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				63297 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				63319 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				63405 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				63410 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				63415 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				63427 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				63454 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				63627 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				63641 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				63655 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				63706 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				63709 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				63788 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				63810 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				63845 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				63852 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				63892 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				63948 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				63949 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				64028 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				64141 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				64166 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				64194 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				64221 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				64245 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				64263 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				64271 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				64300 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				64320 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				64322 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				64341 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				64386 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				64400 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				64419 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				64448 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				64478 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				64483 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				64496 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				64657 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				64665 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				64666 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				64691 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				64723 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				64786 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				64808 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				64902 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				65148 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				65221 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				65226 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				65274 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				65276 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				65278 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				65332 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				65372 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				65401 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				65435 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				65444 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),

                                OTHERS => STD_LOGIC_VECTOR(to_unsigned(2, 8))
                            );
                    
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
                ASSERT (mem_we = '1' OR mem_we = '0') REPORT "o_mem_we in an unexpected state" SEVERITY failure;
            END IF;
            ASSERT (enable_wire = '1' OR enable_wire = '0') REPORT "o_mem_en in an unexpected state" SEVERITY failure;
        END IF;
    END PROCESS;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    createScenario : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '0' THEN
            tb_rst <= scenario_rst(0);
            tb_w <= scenario_w(0);
            tb_start <= scenario_start(0);
            scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_done = '0' REPORT "TEST FALLITO (postreset DONE != 0 )" SEVERITY failure;
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(2, 8)) severity failure; --110001011011:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(2, 8)) severity failure; --110101111000101:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1111001101101111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(2, 8)) severity failure; --0110100101100001:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --011001000001111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1100011110000111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1100111111111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1000010011011:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(2, 8)) severity failure; --01101001101111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8)) severity failure; --101110111100101:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --111100110001101:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1101101001000111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --000001:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --0011011101:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(2, 8)) severity failure; --100110100100111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(2, 8)) severity failure; --110101100101101:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1011000001110001:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(2, 8)) severity failure; --10010100101001:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8)) severity failure; --0100111100011101:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1101001101111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1000001011001:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8)) severity failure; --011011110110111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --01010001010001:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8)) severity failure; --010001100001001:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --010000100000011:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1110011101010101:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --0001011001111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1001000111010011:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(2, 8)) severity failure; --000100000100101:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8)) severity failure; --111111110011001:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(2, 8)) severity failure; --0011001100010111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1010001010111111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1101111111111011:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8)) severity failure; --11110111110101:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8)) severity failure; --0000000001110101:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(2, 8)) severity failure; --0001100101101001:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(2, 8)) severity failure; --011010110111011:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --111000011010111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(2, 8)) severity failure; --100101010110001:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --1110111011111111:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(2, 8)) severity failure; --0010101101111001:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8)) severity failure; --0001001101111011:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(2, 8)) severity failure; --00011101111101:2
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 

        ASSERT false REPORT "Simulation Ended! TEST PASSATO (EXAMPLE)" SEVERITY failure;
    END PROCESS testRoutine;

END projecttb;