LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 1072; 
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00110" & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000" & "11111111111111111000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000000000111111111111111111000000000000000001111111111111111100000000000000000000000000111111111111111111000000001111111111111000000000000000000000000011111111111111111000000000001111111111111111100000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000000001111111111111110000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000000000011111111111111111100000000000000000000000000111111111111111110000000000000000000111111111111111110000000000000011111111111111110000000000000000000000000011111111111111111100000000000000111111111111110000000001111111111110000000011111111111111111000011111111111111111000000000000000000000011111111111111111100000000000000000000000000111111111111111110000000111111111111111111000000000000000000011111111111111100000000000000";
    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000" & "01100010100111101000000000000000001110101010101000100000000000000000000000000011111000111110000000000000000000000000000111110011101101111000000000000000001111110001110001100000000000000000000000000011101000000110001000000000100100110111000000000000000000000000010000110000101011000000000001100100011001011100000000010111100111111001100000000000000000000000000101010100110011110000000000000000000000000001110000001000111000000000000001111011110011100010000000000000000000000000010110010101101001100000000000000000000000000000001101100010010000000000000000000001001011100101111000000000000000000000011001000000100001100000000000000000000000000000000000011110110001100000000000000000000000000100110100111010110000000000000000000000001100111101010000000000000011100111101101010000000000000000000000000011001000000100111100000000000000111100110000110000000001010110010010000000000111011000001001000011110110011000001000000000000000000000010111110001011011100000000000000000000000000010111110100111110000000010011011000001111000000000000000000011110100111010100000000000000";

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (  
				181 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				312 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				349 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				386 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				405 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				419 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				443 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				512 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				581 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				741 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				827 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				984 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				1132 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				1153 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				1168 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				1256 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				1294 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				1487 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				1510 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				1687 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				1699 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				1732 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				1782 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				1952 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				1972 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				1973 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				2008 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				2042 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				2159 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				2218 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				2266 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				2395 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				2574 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				2661 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				2752 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				2820 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				2831 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				2849 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				2938 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				3009 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				3129 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				3140 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				3158 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				3190 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				3240 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				3293 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				3300 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				3353 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				3433 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				3537 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				3595 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				3610 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				3616 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				3731 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				3775 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				3861 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				4033 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				4102 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				4357 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				4425 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				4486 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				4499 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				4511 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				4645 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				4707 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				4719 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				4804 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				4838 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				4911 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				4923 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				5148 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				5203 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				5222 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				5280 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				5281 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				5364 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				5380 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				5475 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				5483 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				5486 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				5567 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				5613 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				5655 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				5661 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				5663 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				5899 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				5905 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				5987 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				6129 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				6186 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				6225 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				6287 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				6379 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				6388 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				6505 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				6629 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				6639 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				6673 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				6734 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				6824 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				6849 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				6930 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				6952 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				6992 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				7209 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				7243 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				7455 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				7569 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				7589 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				7595 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				7636 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				7638 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				7685 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				7714 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				7852 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				7857 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				7887 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				7950 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				8020 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				8052 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				8122 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				8144 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				8168 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				8188 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				8298 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				8593 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				8612 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				8613 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				8757 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				8773 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				8985 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				9029 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				9044 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				9063 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				9129 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				9142 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				9163 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				9314 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				9320 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				9491 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				9617 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				9756 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				9791 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				9821 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				9889 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				9927 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				10068 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				10124 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				10155 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				10195 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				10470 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				10482 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				10518 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				10539 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				10545 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				10604 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				10715 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				10804 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				10950 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				11166 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				11308 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				11435 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				11480 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				11512 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				11522 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				11524 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				11531 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				11545 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				11673 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				11708 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				11730 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				11829 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				11830 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				11855 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				11873 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				11888 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				12004 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				12234 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				12380 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				12421 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				12507 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				12670 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				12923 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				12959 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				12962 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				12965 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				13096 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				13122 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				13181 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				13223 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				13232 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				13279 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				13295 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				13383 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				13384 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				13395 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				13414 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				13480 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				13523 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				13600 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				13614 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				13624 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				13717 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				13854 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				13888 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				13952 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				14022 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				14132 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				14218 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				14331 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				14394 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				14429 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				14450 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				14470 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				14478 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				14586 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				14655 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				14728 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				14771 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				15088 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				15090 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				15211 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				15227 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				15349 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				15398 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				15411 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				15449 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				15467 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				15473 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				15476 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				15593 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				15632 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				15765 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				15802 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				15829 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				16062 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				16317 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				16461 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				16530 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				16532 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				16539 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				16622 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				16677 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				16685 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				16803 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				16814 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				17035 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				17144 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				17428 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				17463 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				17578 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				17586 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				17762 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				17763 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				17766 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				17829 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				17912 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				17925 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				17953 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				17996 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				18129 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				18146 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				18192 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				18239 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				18250 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				18283 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				18363 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				18366 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				18629 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				18659 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				18799 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				18848 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				18910 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				18954 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				19016 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				19150 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				19180 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				19592 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				19637 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				19690 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				19857 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				20004 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				20035 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				20043 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				20080 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				20229 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				20272 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				20364 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				20436 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				20477 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				20479 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				20594 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				20622 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				20831 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				20843 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				20892 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				20898 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				20926 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				21093 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				21138 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				21248 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				21273 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				21340 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				21394 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				21439 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				21454 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				21536 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				21563 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				21565 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				21572 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				21582 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				21642 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				21689 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				21702 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				21719 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				21911 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				21962 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				22005 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				22051 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				22098 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				22148 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				22264 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				22425 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				22443 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				22468 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				22504 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				22533 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				22614 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				22721 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				22722 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				22769 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				22817 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				22861 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				22973 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				22975 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				23027 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				23125 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				23158 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				23379 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				23487 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				23492 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				23517 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				23652 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				23688 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				23699 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				23706 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				23715 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				23745 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				23780 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				23785 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				23807 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				23808 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				23820 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				23873 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				23880 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				23884 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				23925 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				23959 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				24038 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				24065 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				24111 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				24235 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				24326 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				24335 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				24344 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				24430 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				24511 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				24583 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				24624 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				24635 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				24666 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				24769 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				24856 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				24914 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				24932 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				24983 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				25018 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				25110 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				25221 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				25354 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				25628 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				25654 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				25658 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				25668 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				25764 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				25815 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				25909 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				26044 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				26046 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				26049 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				26148 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				26153 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				26159 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				26320 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				26354 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				26577 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				26582 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				26671 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				26722 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				26749 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				26801 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				26816 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				26894 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				27064 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				27108 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				27182 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				27217 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				27244 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				27261 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				27304 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				27466 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				27531 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				27601 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				27777 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				27794 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				27911 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				27947 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				28009 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				28022 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				28038 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				28063 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				28162 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				28163 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				28308 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				28477 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				28569 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				28613 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				28743 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				28748 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				28799 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				28828 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				28885 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				28888 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				28889 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				28901 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				28908 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				28930 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				28931 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				28936 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				28980 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				29030 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				29061 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				29082 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				29118 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				29156 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				29166 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				29314 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				29542 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				29647 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				29688 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				29707 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				29887 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				29944 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				29959 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				30010 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				30043 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				30047 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				30055 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				30092 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				30134 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				30246 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				30380 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				30388 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				30442 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				30576 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				30631 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				30742 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				30750 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				30758 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				30903 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				31062 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				31068 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				31097 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				31139 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				31159 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				31177 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				31211 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				31227 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				31244 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				31252 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				31255 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				31296 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				31372 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				31405 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				31425 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				31489 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				31518 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				31605 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				31670 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				31775 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				31865 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				31910 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				32010 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				32141 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				32283 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				32556 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				32574 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				33131 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				33179 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				33180 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				33245 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				33265 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				33312 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				33343 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				33434 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				33448 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				33479 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				33530 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				33731 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				33765 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				33778 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				33805 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				33897 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				33963 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				33997 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				34282 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				34308 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				34339 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				34378 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				34397 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				34411 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				34430 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				34435 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				34480 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				34483 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				34559 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				34578 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				34720 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				34802 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				34861 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				34877 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				35176 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				35214 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				35307 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				35340 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				35382 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				35443 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				35538 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				35543 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				35794 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				35867 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				35877 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				35912 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				35971 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				36020 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				36199 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				36320 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				36328 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				36342 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				36350 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				36477 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				36599 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				36699 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				36795 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				36852 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				36854 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				36898 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				36937 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				37134 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				37338 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				37402 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				37493 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				37569 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				37608 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				37699 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				37727 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				37789 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				37798 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				37801 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				37812 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				37883 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				37903 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				37956 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				38075 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				38136 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				38178 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				38180 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				38223 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				38329 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				38362 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				38491 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				38533 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				38594 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				38659 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				38753 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				38789 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				38857 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				38876 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				38915 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				39060 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				39074 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				39113 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				39122 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				39295 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				39324 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				39367 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				39371 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				39442 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				39474 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				39496 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				39517 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				39611 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				39625 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				39639 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				39809 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				39810 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				39846 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				39848 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				39853 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				39885 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				39907 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				39998 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				40040 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				40091 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				40095 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				40116 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				40156 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				40163 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				40241 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				40245 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				40261 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				40348 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				40465 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				40546 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				40554 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				40839 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				40844 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				40910 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				40927 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				40953 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				41065 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				41102 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				41126 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				41182 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				41210 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				41251 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				41274 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				41355 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				41379 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				41444 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				41561 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				41573 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				41706 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				41831 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				41929 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				41933 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				42004 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				42033 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				42043 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				42067 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				42095 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				42179 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				42200 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				42269 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				42360 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				42369 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				42461 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				42546 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				42565 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				42604 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				42682 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				42719 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				42767 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				42792 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				42806 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				42862 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				42874 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				42880 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				43064 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				43149 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				43200 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				43456 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				43616 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				43637 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				43835 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				43837 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				43872 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				43959 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				44063 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				44166 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				44222 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				44334 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				44406 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				44407 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				44476 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				44614 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				44619 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				44629 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				44694 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				44696 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				44842 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				44930 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				44977 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				44978 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				45037 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				45091 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				45167 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				45187 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				45251 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				45465 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				45614 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				45695 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				45826 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				45844 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				46027 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				46044 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				46066 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				46085 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				46119 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				46216 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				46276 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				46340 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				46348 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				46454 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				46638 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				46718 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				46840 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				46881 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				46922 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				46940 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				46981 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				46995 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				46996 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				47009 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				47014 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				47025 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				47038 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				47057 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				47129 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				47184 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				47417 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				47476 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				47535 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				47691 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				47714 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				47717 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				47719 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				47780 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				47850 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				47919 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				47958 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				47971 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				48085 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				48167 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				48311 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				48433 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				48511 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				48654 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				48806 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				48818 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				48842 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				48887 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				48888 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				48942 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				48980 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				48986 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				49086 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				49104 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				49123 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				49234 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				49282 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				49354 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				49450 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				49474 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				49534 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				49619 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				49768 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				50022 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				50023 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				50100 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				50129 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				50140 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				50172 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				50239 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				50309 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				50397 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				50520 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				50570 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				50579 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				50626 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				50694 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				50818 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				50865 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				50876 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				50883 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				50892 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				50897 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				50973 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				50997 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				51108 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				51120 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				51145 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				51171 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				51332 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				51383 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				51466 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				51485 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				51518 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				51524 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				51572 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				51580 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				51583 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				51787 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				51843 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				51958 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				52076 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				52198 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				52263 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				52303 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				52310 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				52320 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				52336 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				52395 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				52473 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				52505 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				52562 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				52564 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				52567 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				52580 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				52668 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				52709 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				52711 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				52765 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				52777 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				52806 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				52891 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				52907 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				52910 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				52939 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				52940 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				53049 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				53254 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				53373 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				53393 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				53444 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				53606 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				53610 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				53638 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				53663 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				53743 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				53749 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				53813 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				53864 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				53882 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				53914 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				53966 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				53976 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				54272 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				54287 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				54324 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				54366 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				54459 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				54472 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				54485 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				54527 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				54588 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				54594 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				54607 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				54675 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				54755 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				54762 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				54780 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				54842 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				54850 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				54861 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				54889 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				54983 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				55230 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				55411 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				55529 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				55633 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				55798 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				55894 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				55956 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				55998 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				56063 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				56083 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				56130 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				56140 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				56170 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				56198 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				56217 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				56373 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				56437 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				56487 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				56646 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				56671 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				56757 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				56854 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				56972 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				57060 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				57121 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				57193 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				57284 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				57311 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				57362 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				57392 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				57413 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				57479 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				57508 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				57574 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				57612 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				57647 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				57687 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				57744 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				58019 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				58083 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				58155 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				58506 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				58535 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				58577 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				58612 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				58680 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				58693 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				58719 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				58747 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				58777 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				58789 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				58891 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				58944 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				58964 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				59037 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				59068 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				59077 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				59147 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				59215 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				59254 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				59272 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				59297 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				59341 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				59346 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				59534 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				59633 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				59634 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				59635 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				59696 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				59938 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				60001 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				60076 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				60283 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				60401 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				60563 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				60586 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				60616 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				60629 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				60716 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				60744 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				60808 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				60813 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				60822 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				60910 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				60912 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				61008 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				61051 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				61058 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				61121 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				61168 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				61283 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				61298 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				61480 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				61542 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				61546 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				61589 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				61671 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				61857 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				61910 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				61960 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				62007 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				62033 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				62170 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				62295 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				62439 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				62467 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				62469 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				62518 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				62525 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				62568 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				62628 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				62691 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				62814 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				62849 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				62965 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				63023 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				63032 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				63042 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				63053 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				63061 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				63096 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				63129 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				63187 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				63239 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				63241 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				63310 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				63610 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				63640 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				63689 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				63849 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				63957 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				64010 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				64086 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				64105 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				64123 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				64127 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				64204 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				64336 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				64380 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				64396 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				64426 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				64474 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				64491 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				64892 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				64897 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				64976 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				65084 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				65142 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				65404 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				65467 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),

                                OTHERS => STD_LOGIC_VECTOR(to_unsigned(183, 8))
                            );
                    
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
                ASSERT (mem_we = '1' OR mem_we = '0') REPORT "o_mem_we in an unexpected state" SEVERITY failure;
            END IF;
            ASSERT (enable_wire = '1' OR enable_wire = '0') REPORT "o_mem_en in an unexpected state" SEVERITY failure;
        END IF;
    END PROCESS;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    createScenario : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '0' THEN
            tb_rst <= scenario_rst(0);
            tb_w <= scenario_w(0);
            tb_start <= scenario_start(0);
            scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_done = '0' REPORT "TEST FALLITO (postreset DONE != 0 )" SEVERITY failure;
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 100010100111101:183 -> 01 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 1101010101010001:183 -> 01 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 01111100011111:183 -> 00 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 1110011101101111:183 -> 11 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 111100011100011:183 -> 11 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 1101000000110001:183 -> 01 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 00100110111:183 -> 01 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 000110000101011:183 -> 10 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 001000110010111:183 -> 11 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 1111001111110011:183 -> 10 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 0101010011001111:183 -> 01 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 1110000001000111:183 -> 00 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 1101111001110001:183 -> 11 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 1100101011010011:183 -> 10 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 0110110001001:183 -> 00 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 1001011100101111:183 -> 00 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 0010000001000011:183 -> 11 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 0000111101100011:183 -> 00 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 011010011101011:183 -> 10 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 000110011110101:183 -> 00 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 10011110110101:183 -> 11 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 0010000001001111:183 -> 11 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 110011000011:183 -> 11 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 1011001001:183 -> 10 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 111011000001001:183 -> 00 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 110110011000001:183 -> 11 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 1111100010110111:183 -> 10 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 011111010011111:183 -> 01 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 0011011000001111:183 -> 01 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8)) severity failure; -- 1101001110101:183 -> 11 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 

        ASSERT false REPORT "Simulation Ended! TEST PASSATO (EXAMPLE)" SEVERITY failure;
    END PROCESS testRoutine;

END projecttb;