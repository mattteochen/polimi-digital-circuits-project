LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 2914; 
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00110" & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000" & "11111111111111111100000000000000000000000000111111111111111111000000000000000000011111111111111111100000000111111111111111111000000011111111111111111100000000000000111111111111111111000000000111111111111111100000000000000000000000000001111111111111111000000000001111111111111111110000000000000000000000000000011111111111111111100000000000000000000111111111111111111000000000000111111111111111110000000000000000000000000000001111111111111000000000000000000111111111111111110000000000000000000011111111111111111000000000000000011111111111111111000000000000000000000000000111111111111111111000000000111111111100000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000000000111111111111111000000000000000000000000001111111111111111000000000000000000011111111111111111100000000000000011111111111111111100000000000000000000111111111111111111000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000000011111111111110000000000000000111111111111111110000000000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000001111111111111111100000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000011111111111111111000000000000000000111111111111111110000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000000001111111111111100000001111111111111111100000000000000000001111111111111111110000000111111111111111111000000000000011111111111111100000000000001111111111111111100000000000000000000000000000111111111111110000000000000000000001111111111111111110000000000000000000000000001111111111111110000000000000000000000000000001111111111111111110000000000000000000000000000111111111111111000000000000011111111111111111100000000000000000000000000111111111111111111000000000111111111111110000000000000000000011111111111111111100000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000111111111111111100000000000000000111111111111111111000000000000000000011111111111111111100000000000000000111111111111111110000000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000001111111111111111100000000000000011111111111111111000000000000000000111111111111111111000000011111111111111111100000000001111111111111111100000000000000000000000000000011111111111111111000000000000011111111111111111100000000000000000001111111111111111000000000000000000001111111111111111100000000000000011111111111111111000000000011111111111111111100000000000000000000011111111111111111100000000000000001111111111111111100000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000001111111111111111100000000000011111111111111111100000000";
    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000" & "10001010011111100100000000000000000000000000010001011100101011000000000000000000010000000000000100100000000001110110100001001000000010101000100100101100000000000000010110101001101011000000000000111111000110100000000000000000000000000001101010000110001000000000000101100100111101110000000000000000000000000000010101001111000011100000000000000000000101110000111001011000000000000101011001100101110000000000000000000000000000000000001011011000000000000000000110110101001111110000000000000000000000100000000101001000000000000000010001110101001001000000000000000000000000000100111111101000001000000000000110100100000000000000000000101110111011101110000000000000000000000000110010000110110010000000000000000000000000000110110101000101000000000000000000000000000110011010110101000000000000000000000001000111000001100000000000000010000110001110110100000000000000000000110011000101000001000000000000010001110011001010000000000000000000000011110100011000101100000000000000000000000000010111001000110000000000000000011000111110101010000000000000000000000000000000100110111101010110000000000000000000000000010001001001110111100000000000000000001101100101011100100000000000000000000000000011100011001000110100000000000000000000000010011011101011101100000000000000000000000000100100110110100001000000000000001010111000111001000000000000000000101001101000110010000000000000000000100100101111000000000000000000000000000010001100111010000000000000000000000000001011011100101100000001001000010110000100000000000000000000000000100100111010000000101001101110100111000000000000001001100101101100000000000001000011110110001100000000000000000000000000000101011101111110000000000000000000001111100100011101110000000000000000000000000000111000101000010000000000000000000000000000001010100001110111010000000000000000000000000000001011000100001000000000000001001100011110011100000000000000000000000000110001101101101001000000000011101110000010000000000000000000010011010100010111100000000000000000000000010100001000100000000000000000000000010011100001110010000000000000000000000000000110100001101010000000000000000000001011110111100000000000000000110111011000111011000000000000000000010011011011101101100000000000000000100101101010000010000000000000000000000000001010000010011101010000000000000000000000010101101010000111000000000000000000101110001000010100000000000000011101001111001101000000000000000000111101011110010101000000000110100010001010100000000001111000100111011100000000000000000000000000000010001010001110111000000000000001001011011101111100000000000000000000001100110100101000000000000000000000111101111011011100000000000000011110111010001001000000000000110000111101101100000000000000000000011001110011011101100000000000000001111111010101101100000000000000000001101101111010001110000000000000000000000000111011001111111100000000000000000000010011101101110101100000001001100110110111100000000000000100101101100111100000000";

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (  
				1 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				20 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				83 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				176 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				179 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				232 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				337 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				342 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				473 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				529 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				531 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				612 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				614 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				660 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				688 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				712 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				749 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				751 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				810 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				833 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				838 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				877 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				933 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				969 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				1036 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				1052 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				1062 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				1181 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				1184 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				1208 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				1222 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				1279 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				1299 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				1318 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				1425 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				1557 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				1602 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				1614 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				1633 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				1643 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				1836 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				1903 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				1922 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				1997 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				2087 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				2088 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				2100 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				2103 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				2113 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				2163 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				2189 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				2225 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				2245 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				2277 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				2381 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				2470 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				2497 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				2524 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				2607 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				2613 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				2623 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				2761 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				2784 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				2798 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				2887 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				2934 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				2957 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				3026 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				3040 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				3044 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				3062 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				3090 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				3167 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				3297 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				3298 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				3377 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				3395 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				3461 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				3543 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				3577 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				3609 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				3626 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				3744 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				3749 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				3774 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				3786 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				3800 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				3801 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				3830 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				3847 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				3860 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				3874 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				3945 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				3952 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				3982 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				3988 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				4012 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				4013 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				4014 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				4031 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				4064 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				4096 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				4162 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				4195 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				4263 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				4279 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				4302 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				4359 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				4400 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				4507 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				4525 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				4545 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				4702 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				4745 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				4783 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				4953 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				4965 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				5001 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				5021 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				5040 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				5042 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				5156 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				5180 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				5268 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				5269 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				5352 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				5390 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				5441 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				5515 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				5516 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				5573 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				5600 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				5627 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				5664 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				5780 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				5916 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				5924 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				6042 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				6052 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				6070 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				6137 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				6174 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				6205 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				6220 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				6252 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				6300 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				6329 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				6378 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				6401 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				6405 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				6412 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				6556 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				6565 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				6617 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				6685 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				6731 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				6746 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				6748 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				6778 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				6796 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				6806 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				6832 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				6894 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				6941 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				6949 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				6985 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				7059 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				7068 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				7200 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				7204 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				7277 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				7301 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				7307 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				7320 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				7326 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				7374 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				7384 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				7429 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				7440 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				7481 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				7535 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				7694 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				7699 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				7704 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				7733 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				7744 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				7773 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				7795 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				7816 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				7861 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				7886 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				8018 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				8036 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				8040 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				8149 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				8151 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				8227 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				8278 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				8317 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				8424 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				8437 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				8446 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				8501 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				8503 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				8559 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				8609 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				8626 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				8678 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				8755 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				8896 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				8928 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				9038 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				9075 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				9125 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				9127 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				9169 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				9173 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				9176 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				9201 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				9216 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				9297 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				9329 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				9390 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				9398 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				9444 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				9446 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				9461 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				9529 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				9546 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				9574 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				9650 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				9685 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				9696 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				9801 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				9862 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				9867 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				9892 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				9920 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				10043 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				10046 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				10116 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				10120 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				10130 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				10161 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				10189 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				10218 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				10232 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				10266 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				10273 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				10275 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				10381 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				10401 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				10429 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				10489 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				10493 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				10516 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				10530 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				10532 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				10575 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				10599 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				10622 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				10684 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				10729 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				10758 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				10779 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				10885 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				10904 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				11037 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				11065 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				11081 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				11150 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				11197 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				11206 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				11239 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				11242 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				11294 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				11302 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				11308 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				11706 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				11727 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				11736 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				11792 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				11844 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				11997 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				12006 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				12111 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				12141 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				12143 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				12155 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				12163 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				12205 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				12316 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				12394 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				12395 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				12424 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				12461 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				12508 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				12513 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				12536 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				12592 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				12672 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				12696 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				12710 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				12808 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				12873 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				12888 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				12902 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				12964 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				12985 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				13008 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				13074 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				13079 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				13094 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				13095 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				13102 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				13120 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				13309 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				13313 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				13408 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				13506 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				13528 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				13587 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				13592 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				13613 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				13645 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				13728 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				13743 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				13818 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				13868 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				13870 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				13873 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				13929 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				13937 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				13974 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				14019 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				14033 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				14073 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				14088 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				14101 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				14122 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				14226 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				14240 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				14247 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				14251 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				14263 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				14285 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				14292 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				14329 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				14381 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				14410 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				14467 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				14534 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				14580 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				14584 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				14706 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				14731 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				14808 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				14820 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				14907 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				14938 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				14963 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				15056 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				15134 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				15190 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				15254 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				15260 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				15389 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				15514 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				15521 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				15579 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				15610 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				15651 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				15701 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				15758 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				15780 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				15798 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				15849 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				15916 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				15922 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				15944 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				16019 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				16030 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				16235 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				16249 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				16284 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				16335 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				16401 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				16447 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				16459 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				16482 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				16532 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				16547 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				16548 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				16569 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				16597 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				16718 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				16770 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				16787 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				16849 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				16863 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				16898 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				16982 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				17007 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				17014 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				17087 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				17094 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				17156 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				17457 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				17615 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				17639 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				17646 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				17665 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				17710 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				17714 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				17744 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				17831 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				17903 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				18014 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				18108 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				18233 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				18234 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				18241 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				18266 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				18335 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				18465 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				18569 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				18620 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				18649 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				18666 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				18739 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				18742 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				18743 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				18796 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				18831 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				18867 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				18875 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				18967 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				19008 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				19063 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				19164 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				19250 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				19264 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				19385 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				19388 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				19390 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				19398 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				19430 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				19443 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				19457 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				19481 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				19498 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				19511 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				19514 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				19515 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				19532 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				19577 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				19592 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				19657 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				19664 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				19672 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				19712 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				19720 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				19748 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				19837 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				19859 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				19941 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				19956 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				19984 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				19989 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				19997 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				20034 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				20046 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				20049 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				20054 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				20105 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				20125 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				20126 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				20145 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				20307 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				20314 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				20345 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				20370 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				20373 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				20374 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				20397 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				20505 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				20524 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				20627 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				20821 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				20832 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				20858 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				20903 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				20939 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				21084 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				21106 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				21161 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				21182 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				21194 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				21225 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				21285 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				21330 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				21400 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				21407 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				21414 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				21421 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				21468 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				21551 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				21572 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				21597 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				21635 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				21666 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				21741 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				21754 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				21770 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				21774 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				21815 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				21874 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				21892 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				21928 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				21929 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				21966 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				22067 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				22146 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				22236 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				22257 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				22265 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				22356 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				22439 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				22441 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				22522 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				22753 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				22810 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				22813 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				22831 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				22905 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				22939 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				22969 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				23188 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				23214 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				23216 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				23337 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				23360 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				23406 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				23480 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				23550 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				23602 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				23661 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				23673 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				23681 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				23831 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				23857 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				23902 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				23922 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				23923 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				23994 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				23996 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				24021 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				24060 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				24074 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				24157 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				24208 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				24324 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				24378 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				24389 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				24452 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				24456 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				24529 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				24542 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				24582 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				24602 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				24651 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				24657 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				24751 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				24773 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				24878 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				24915 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				24919 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				24923 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				25066 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				25244 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				25280 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				25367 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				25411 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				25418 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				25442 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				25470 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				25545 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				25611 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				25640 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				25773 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				25815 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				25884 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				25933 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				25937 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				25952 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				26014 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				26029 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				26058 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				26086 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				26188 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				26231 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				26253 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				26358 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				26372 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				26418 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				26428 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				26446 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				26451 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				26559 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				26571 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				26617 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				26640 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				26786 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				26852 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				26892 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				26908 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				26915 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				26925 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				26994 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				27005 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				27026 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				27048 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				27062 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				27068 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				27101 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				27117 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				27136 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				27169 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				27185 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				27208 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				27256 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				27297 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				27335 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				27358 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				27389 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				27420 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				27425 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				27430 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				27443 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				27466 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				27503 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				27506 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				27545 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				27583 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				27617 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				27636 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				27647 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				27657 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				27789 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				27841 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				27905 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				27918 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				27985 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				27986 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				27987 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				27992 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				28071 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				28116 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				28217 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				28228 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				28276 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				28290 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				28308 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				28309 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				28334 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				28337 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				28338 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				28401 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				28424 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				28434 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				28438 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				28458 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				28519 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				28543 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				28640 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				28644 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				28694 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				28865 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				28954 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				28992 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				29002 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				29089 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				29138 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				29194 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				29228 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				29229 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				29238 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				29269 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				29352 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				29437 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				29500 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				29580 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				29595 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				29647 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				29675 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				29746 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				29905 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				29973 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				29994 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				30000 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				30016 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				30037 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				30071 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				30107 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				30151 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				30165 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				30218 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				30229 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				30314 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				30347 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				30387 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				30407 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				30432 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				30450 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				30452 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				30461 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				30469 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				30483 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				30496 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				30523 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				30563 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				30564 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				30614 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				30737 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				30742 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				30751 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				30818 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				30942 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				30973 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				30981 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				31017 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				31046 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				31052 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				31098 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				31111 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				31176 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				31206 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				31257 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				31273 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				31358 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				31377 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				31408 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				31460 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				31566 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				31577 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				31607 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				31614 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				31681 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				31723 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				31769 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				31827 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				31929 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				31948 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				31961 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				31964 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				32044 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				32064 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				32090 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				32160 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				32190 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				32217 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				32235 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				32238 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				32252 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				32303 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				32366 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				32453 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				32468 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				32488 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				32626 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				32667 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				32676 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				32785 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				32830 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				32834 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				32900 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				32916 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				32969 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				32994 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				33115 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				33151 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				33156 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				33160 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				33164 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				33202 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				33230 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				33394 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				33437 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				33456 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				33499 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				33509 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				33528 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				33554 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				33556 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				33567 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				33571 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				33587 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				33613 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				33658 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				33718 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				33763 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				33778 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				33815 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				33839 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				33870 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				33950 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				33969 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				33970 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				33990 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				34048 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				34071 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				34079 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				34137 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				34138 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				34161 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				34176 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				34225 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				34262 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				34335 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				34348 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				34489 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				34530 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				34541 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				34690 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				34777 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				34801 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				34838 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				34951 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				34967 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				34999 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				35012 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				35054 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				35100 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				35134 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				35159 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				35163 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				35200 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				35244 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				35276 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				35323 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				35425 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				35480 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				35482 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				35538 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				35580 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				35587 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				35596 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				35619 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				35641 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				35723 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				35787 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				35806 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				35866 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				35882 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				35908 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				35930 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				35954 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				35966 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				36005 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				36012 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				36065 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				36171 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				36201 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				36235 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				36285 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				36296 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				36333 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				36340 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				36524 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				36534 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				36547 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				36614 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				36707 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				36712 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				36725 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				36728 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				36742 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				36782 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				36853 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				36915 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				36960 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				36984 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				37058 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				37115 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				37187 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				37266 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				37305 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				37332 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				37402 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				37425 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				37468 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				37565 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				37623 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				37650 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				37659 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				37722 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				37904 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				38035 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				38037 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				38081 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				38118 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				38150 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				38157 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				38180 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				38182 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				38187 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				38196 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				38267 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				38283 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				38348 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				38376 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				38381 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				38385 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				38417 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				38518 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				38576 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				38583 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				38660 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				38695 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				38734 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				38765 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				38769 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				38774 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				38799 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				38801 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				38806 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				38850 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				38863 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				38951 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				39012 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				39051 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				39056 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				39077 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				39100 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				39130 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				39143 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				39233 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				39272 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				39283 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				39296 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				39337 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				39356 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				39371 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				39375 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				39399 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				39501 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				39520 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				39522 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				39674 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				39726 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				39771 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				39799 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				39818 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				39826 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				39876 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				39912 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				39915 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				39927 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				39977 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				40013 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				40017 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				40049 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				40224 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				40227 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				40255 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				40259 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				40303 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				40321 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				40323 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				40354 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				40442 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				40478 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				40554 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				40576 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				40683 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				40729 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				40751 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				40763 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				40773 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				40809 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				40864 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				40870 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				40879 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				40881 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				40915 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				40982 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				41000 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				41052 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				41119 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				41165 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				41183 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				41221 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				41268 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				41310 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				41380 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				41394 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				41421 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				41479 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				41522 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				41524 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				41546 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				41575 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				41675 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				41712 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				41863 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				41905 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				41943 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				42008 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				42019 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				42037 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				42212 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				42260 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				42267 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				42276 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				42345 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				42442 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				42474 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				42506 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				42556 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				42592 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				42605 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				42630 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				42652 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				42659 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				42675 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				42716 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				42747 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				42752 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				42765 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				42783 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				42814 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				42862 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				42877 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				42940 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				42988 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				42996 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				43006 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				43018 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				43031 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				43066 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				43099 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				43118 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				43147 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				43199 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				43523 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				43551 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				43586 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				43591 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				43593 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				43599 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				43722 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				43798 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				43808 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				43860 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				43898 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				43901 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				43908 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				43917 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				43950 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				43982 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				43996 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				44016 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				44082 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				44091 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				44095 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				44144 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				44176 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				44235 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				44382 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				44415 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				44417 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				44455 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				44514 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				44519 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				44560 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				44583 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				44585 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				44605 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				44631 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				44797 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				44817 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				44839 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				45014 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				45060 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				45095 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				45156 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				45162 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				45167 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				45185 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				45194 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				45205 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				45221 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				45265 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				45371 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				45374 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				45394 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				45396 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				45424 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				45442 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				45447 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				45470 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				45475 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				45517 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				45556 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				45584 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				45596 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				45616 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				45651 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				45655 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				45656 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				45712 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				45776 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				45802 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				45859 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				45881 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				45896 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				45911 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				46020 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				46054 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				46071 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				46122 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				46150 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				46314 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				46315 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				46437 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				46453 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				46652 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				46667 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				46753 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				46782 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				46807 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				46952 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				46965 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				46981 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				46995 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				47004 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				47115 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				47141 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				47169 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				47174 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				47184 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				47192 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				47195 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				47311 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				47380 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				47398 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				47430 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				47489 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				47587 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				47632 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				47689 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				47754 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				47903 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				47967 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				47997 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				48027 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				48230 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				48299 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				48370 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				48402 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				48435 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				48497 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				48511 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				48520 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				48556 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				48588 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				48749 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				48750 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				48768 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				48822 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				48860 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				48884 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				48911 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				48930 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				48948 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				48992 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				49050 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				49121 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				49203 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				49240 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				49300 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				49312 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				49320 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				49335 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				49364 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				49473 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				49502 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				49538 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				49557 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				49621 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				49636 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				49714 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				49729 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				49865 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				49867 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				49882 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				49916 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				49920 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				49970 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				49982 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				49997 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				50026 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				50059 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				50097 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				50213 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				50220 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				50249 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				50259 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				50260 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				50300 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				50321 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				50387 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				50415 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				50483 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				50490 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				50512 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				50526 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				50553 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				50588 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				50594 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				50601 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				50606 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				50624 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				50632 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				50718 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				50739 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				50740 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				50954 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				51028 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				51129 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				51179 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				51192 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				51219 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				51220 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				51226 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				51264 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				51267 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				51272 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				51310 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				51351 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				51372 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				51437 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				51479 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				51613 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				51637 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				51698 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				51718 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				51754 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				51780 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				51796 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				51803 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				51921 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				51924 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				51946 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				52044 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				52074 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				52153 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				52173 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				52186 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				52245 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				52328 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				52344 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				52461 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				52462 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				52511 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				52543 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				52562 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				52641 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				52668 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				52712 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				52746 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				52761 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				52780 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				52842 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				52906 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				52966 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				53036 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				53098 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				53137 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				53210 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				53211 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				53312 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				53356 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				53372 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				53390 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				53408 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				53469 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				53498 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				53532 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				53589 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				53625 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				53780 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				53821 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				53882 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				54021 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				54110 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				54111 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				54155 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				54167 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				54168 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				54274 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				54299 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				54336 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				54388 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				54390 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				54442 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				54449 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				54461 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				54483 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				54538 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				54548 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				54612 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				54613 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				54738 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				54780 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				54870 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				55065 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				55270 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				55274 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				55563 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				55584 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				55594 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				55623 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				55750 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				55782 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				55786 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				55794 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				55905 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				55943 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				55983 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				55997 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				56067 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				56123 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				56169 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				56182 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				56185 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				56273 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				56342 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				56347 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				56387 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				56431 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				56478 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				56502 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				56644 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				56655 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				56691 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				56695 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				56697 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				56708 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				56737 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				56777 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				56792 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				56854 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				56954 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				57001 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				57003 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				57058 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				57093 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				57160 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				57169 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				57228 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				57349 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				57396 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				57407 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				57414 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				57416 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				57421 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				57442 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				57460 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				57518 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				57526 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				57626 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				57692 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				57756 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				57759 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				57867 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				57882 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				57905 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				57911 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				57982 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				58039 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				58087 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				58095 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				58145 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				58199 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				58323 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				58348 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				58355 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				58380 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				58400 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				58516 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				58542 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				58552 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				58596 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				58647 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				58754 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				58829 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				58881 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				58915 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				58916 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				58919 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				58942 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				59168 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				59185 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				59215 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				59240 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				59251 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				59346 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				59415 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				59420 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				59476 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				59602 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				59623 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				59659 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				59773 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				59802 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				59871 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				59900 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				59917 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				59919 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				59953 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				60001 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				60007 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				60163 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				60334 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				60350 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				60376 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				60379 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				60453 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				60497 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				60558 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				60578 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				60587 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				60604 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				60693 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				60769 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				60786 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				60802 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				60852 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				60893 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				60901 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				60970 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				60994 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				61004 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				61016 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				61053 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				61152 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				61213 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				61257 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				61265 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				61319 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				61360 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				61379 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				61383 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				61416 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				61434 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				61499 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				61514 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				61565 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				61566 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				61568 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				61614 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				61644 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				61659 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				61663 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				61755 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				61779 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				61789 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				61848 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				61896 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				61904 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				61945 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				61960 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				61973 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				62040 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				62066 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				62166 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				62213 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				62265 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				62269 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				62316 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				62325 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				62403 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				62405 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				62565 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				62594 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				62642 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				62671 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				62704 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				62738 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				62892 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				62932 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				62942 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				63042 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				63098 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				63107 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				63111 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				63129 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				63147 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				63209 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				63249 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				63286 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				63294 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				63323 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				63334 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				63341 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				63410 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				63425 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				63452 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				63482 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				63567 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				63635 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				63646 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				63706 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				63713 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				63719 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				63735 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				63794 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				63822 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				63874 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				63881 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				63883 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				63985 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				64029 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				64036 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				64083 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				64095 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				64179 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				64202 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				64242 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				64257 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				64270 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				64289 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				64354 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				64369 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				64467 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				64508 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				64519 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				64569 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				64634 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				64711 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				64789 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				64833 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				64835 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				64893 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				64910 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				64965 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				65025 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				65087 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				65151 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				65160 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				65179 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				65206 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				65251 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				65353 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				65424 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				65426 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				65436 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				65477 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				65531 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),

                                OTHERS => STD_LOGIC_VECTOR(to_unsigned(207, 8))
                            );
                    
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
                ASSERT (mem_we = '1' OR mem_we = '0') REPORT "o_mem_we in an unexpected state" SEVERITY failure;
            END IF;
            ASSERT (enable_wire = '1' OR enable_wire = '0') REPORT "o_mem_en in an unexpected state" SEVERITY failure;
        END IF;
    END PROCESS;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    createScenario : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '0' THEN
            tb_rst <= scenario_rst(0);
            tb_w <= scenario_w(0);
            tb_start <= scenario_start(0);
            scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_done = '0' REPORT "TEST FALLITO (postreset DONE != 0 )" SEVERITY failure;
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0010100111111001:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0001011100101011:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0000000000001001:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1110110100001001:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1010001001001011:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(166, 8)) severity failure; -- 0110101001101011:166->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 01111110001101:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(166, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 01010000110001:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0110010011110111:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1010011110000111:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1110000111001011:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 101100110010111:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 00001011011:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 011010100111111:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 100000000101001:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 001110101001001:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0111111101000001:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 01101001:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 111011101110111:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 001000011011001:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0110101000101:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 10011010110101:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0010001110000011:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0001100011101101:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0011000101000001:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 00111001100101:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1101000110001011:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 11100100011:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 100011111010101:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0011011110101011:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0010010011101111:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 011001010111001:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1000110010001101:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0110111010111011:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0100110110100001:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 010111000111001:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 100110100011001:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 000100100101111:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 001000110011101:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 110111001011:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 010000101100001:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0000010010011101:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1001101110100111:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0011001011011:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 000111101100011:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 101110111111:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1110010001110111:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1100010100001:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1010000111011101:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1011000100001:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0011000111100111:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0001101101101001:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 110111000001:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0110101000101111:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 000101000010001:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 001110000111001:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0011010000110101:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 00010111101111:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0111011000111011:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0110110111011011:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 010110101000001:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1000001001110101:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0101101010000111:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 011100010000101:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 101001111001101:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1101011110010101:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8)) severity failure; -- 1101000100010101:72->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 110001001110111:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 001010001110111:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0010110111011111:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 01100110100101:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 111011110110111:207->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 110111010001001:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1100001111011011:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0011100110111011:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 111110101011011:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0110111101000111:207->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1110110011111111:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 0111011011101011:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 011001101101111:207->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- 1001011011001111:207->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 

        ASSERT false REPORT "Simulation Ended! TEST PASSATO (EXAMPLE)" SEVERITY failure;
    END PROCESS testRoutine;

END projecttb;