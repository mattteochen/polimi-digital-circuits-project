LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 3363; 
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00110" & "0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000" & "1111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000111111111111111111000000000000000000000111111111111111110000000000011111111111111110000000000000000000111111111111111111000000000000000000000000111111111111111000000000000011111111111111100000000000000000000000111111111111111000000000000000111111111111111110000000000000000000000000000011111111111111111100000000000000000000000000000111111111111111111000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000001111111111111111000000000000000000000000111111111111100000000000000000000011111111111111111100000000000000000000000000000011111111111111111100000000000000000111111111111111111000000011111111111111111100000000000011111111111111111100000000000000000000000001111111111111111110000000001111111111111111100000001111111111111111000000000011111111111111111100000000000000000000000001111111111111111100000000000111111111111111111000000000000111111111111111111000000000000000000111111111111111100000000000000000000000000000111111111111111111000000000111111111111111000000000000111111111111111111000000000000000000000000001111111111111111100000000000000000011111111111111111100000000000111111111111111110000000000000000000111111111111111100000000000000000000000000111111111111111110000000000000000000000000000001111111111111111110000000011111111111111100000000000000001111111111111111110000000001111111111111111110000000000000011111111111111111000000000000000000000001111111111111111110000000000001111111111111111000000001111111111111111110000000111111111111111111000000000000001111111111111111000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000000001111111111111111100000001111111111111111110000000000000000000000000000000111111111111111110000000000000000000000000000011111111111111111100000000000000001111111111111111000000000000111111111111111110000000000000000000000000000111111111111111111000000000000000011111111111111111100000000000011111111111111111100000000000000111111111111111100000000000000000011111111111111111100000001111111111111110000000000000000000000000011111111111111111100000001111111111111000000000000000000000001111111111111111000000000000000000011111111111111111000000000000000000111111111111111111000000000000000000001111111111111111110000000000000001111111111111111110000000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000011111111111111110000000000000000000000000000111111111111111111000000000000000000000000000001111111111111111110000000000011111111111111110000000000001111111111111111110000000000000000001111111111111110000000000111111111111111110000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000111111111111111111000000000000000000000000000000111111111111111100000000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000011111111111111000000000000000000011111111111111110000000111111111111111111000000000000000000000000000000111111111111111111000000000000000000000000000011111111111111111100000000000000000000000000000111111111111110000000000000000000000000000001111111111111110000000000000000000000000000001111111111111111100000000000000000";
    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000" & "0100011100111001110000000000000000000000000000110001000101110000000000000000000000000010100111011011000000000101111110100101111000000000000000000000000001110000000010000000000011011111001000110000000000000000000010001111001000001000000000000000000000000011100101110001000000000000011100010101101100000000000000000000000011011101100011000000000000000000010001101011010000000000000000000000000000010010001010111111100000000000000000000000000000110001001001010101000000000000011100110100011001100000000000000000000000010010110010100010100000000000000000001111111001000011000000000000000000000000111111001001100000000000000000000000010000000000011100000000000000000000000000000011001100111011010100000000000000000101010101001001111000000010001011010101010100000000000001100000111010111100000000000000000000000000100110000001111110000000000000111110011100100000001110000001011101000000000000110101111001110100000000000000000000000000111010000011111100000000000001000100111100101000000000000000110111110011111000000000000000000100100111010011100000000000000000000000000000000100111110110111000000000100101000100111000000000000000101100111111011000000000000000000000000001100111011010100100000000000000000011011111010111001100000000000111011001101101010000000000000000000011000100000111100000000000000000000000000110001101010100110000000000000000000000000000001001111001110100010000000000011110101100100000000000000001100001010011110010000000000100011001111011110000000000000011110011000100111000000000000000000000001111000100010010110000000000001010011001100011000000001100111100101101110000000011000011111010101000000000000001100001100110011000000000101010000000010100000000000000000000000010001001001010011100000000000000000000001000111010111011100000000000000000000000000001000000001000110100000000100111100010111010000000000000000000000000000000001001010010010110000000000000000000000000000011111000110100111100000000000000001111100010111101000000000000101010010110000010000000000000000000000000000001001001011101101000000000000000001000001010010011100000000000010100100110010111100000000000000001101100000010100000000000000000010110000100110000100000000001111000001110000000000000000000000000010010101001010101100000000110000000001000000000000000000000000000000000000011000000000000000000010001000011001001000000000000000000010110110010100111000000000000000000001100010000011010110000000000000001100101000000101110000000000000000000000000001011110001011010100000000000000000000000001001010010010000100000000001110111010111110000000000000000000000000000001111000111000011000000000000000000000000000000001111001011101010000000000001100100101100010000000000000010010010011010110000000000000000001001100111011110000000000111110111011001010000000000000000000000000010011100111011101000000000000000000000001111010101001000110000000000000001000001001110101000000000000000000000000000000000000010101000100000000000000000000000000001000111110001111110000000000000000000000110000111111100110000000000000000000000000010001011011010010000000000000000001001100000011000000000000000000001011010111100110000000111011110001111111000000000000000000000000000000001010100011110111000000000000000000000000000000110101001000101100000000000000000000000000000011010000101110000000000000000000000000000001000110001001010000000000000000000000000000000111110101000100100000000000000000";

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (  
				0 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				11 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				29 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				35 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				39 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				65 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				106 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				165 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				208 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				224 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				229 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				241 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				267 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				279 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				295 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				325 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				352 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				387 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				419 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				462 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				468 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				502 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				541 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				617 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				635 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				643 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				676 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				730 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				742 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				799 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				847 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				869 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				909 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				911 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				941 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				960 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				964 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				986 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				999 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				1048 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				1059 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				1085 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				1225 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				1250 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				1268 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				1335 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				1342 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				1364 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				1533 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				1538 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				1564 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				1575 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				1587 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				1610 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				1758 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				1866 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				1896 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				1898 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				1993 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				2017 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				2035 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				2036 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				2090 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				2103 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				2112 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				2143 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				2146 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				2151 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				2172 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				2214 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				2288 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				2294 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				2299 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				2312 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				2316 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				2466 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				2488 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				2515 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				2534 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				2538 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				2543 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				2616 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				2628 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				2634 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				2668 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				2713 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				2779 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				2821 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				2823 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				2899 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				2976 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				3040 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				3104 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				3227 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				3240 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				3243 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				3343 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				3438 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				3451 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				3489 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				3549 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				3563 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				3652 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				3657 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				3718 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				3738 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				3746 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				3796 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				3848 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				3863 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				3897 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				3921 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				3959 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				4000 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				4038 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				4084 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				4139 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				4142 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				4155 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				4218 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				4220 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				4234 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				4279 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				4336 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				4342 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				4373 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				4394 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				4404 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				4465 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				4534 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				4592 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				4623 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				4627 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				4753 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				4771 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				4772 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				4775 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				4787 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				4840 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				4933 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				4991 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				5003 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				5051 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				5104 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				5169 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				5174 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				5249 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				5282 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				5407 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				5434 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				5447 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				5683 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				5685 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				5701 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				5842 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				5843 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				5902 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				5903 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				5906 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				5915 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				5947 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				5957 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				5970 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				5999 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				6005 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				6085 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				6095 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				6190 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				6230 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				6237 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				6326 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				6329 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				6359 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				6443 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				6490 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				6529 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				6530 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				6581 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				6586 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				6615 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				6654 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				6670 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				6677 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				6692 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				6710 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				6748 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				6806 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				6880 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				6906 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				6947 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				6958 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				7000 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				7054 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				7206 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				7228 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				7255 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				7259 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				7260 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				7287 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				7344 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				7356 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				7417 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				7474 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				7493 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				7504 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				7562 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				7595 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				7599 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				7614 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				7667 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				7752 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				7764 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				7769 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				7790 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				7815 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				7818 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				7870 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				7889 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				7946 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				7952 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				8019 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				8104 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				8136 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				8146 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				8151 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				8186 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				8190 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				8192 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				8238 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				8270 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				8275 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				8294 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				8300 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				8303 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				8319 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				8337 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				8339 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				8400 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				8461 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				8467 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				8470 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				8476 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				8496 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				8508 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				8512 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				8570 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				8578 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				8603 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				8735 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				8739 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				8741 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				8753 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				8772 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				8835 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				8892 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				8918 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				8935 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				9027 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				9040 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				9046 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				9058 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				9075 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				9077 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				9110 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				9146 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				9155 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				9294 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				9342 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				9379 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				9400 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				9422 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				9443 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				9513 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				9526 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				9551 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				9554 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				9581 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				9592 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				9598 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				9695 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				9703 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				9865 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				9875 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				9883 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				9886 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				9899 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				9907 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				9913 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				9933 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				9944 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				9982 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				9986 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				10021 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				10085 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				10136 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				10168 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				10213 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				10251 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				10254 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				10278 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				10345 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				10396 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				10408 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				10671 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				10683 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				10685 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				10738 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				10766 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				10859 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				10867 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				10921 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				11059 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				11084 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				11168 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				11178 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				11221 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				11230 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				11259 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				11399 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				11519 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				11575 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				11678 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				11700 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				11786 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				11811 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				11877 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				11909 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				11970 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				12015 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				12024 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				12057 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				12061 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				12093 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				12118 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				12131 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				12153 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				12178 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				12359 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				12361 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				12368 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				12374 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				12391 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				12400 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				12434 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				12441 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				12453 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				12513 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				12549 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				12595 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				12614 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				12641 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				12648 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				12656 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				12727 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				12765 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				12893 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				12936 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				12976 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				13069 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				13100 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				13120 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				13124 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				13134 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				13173 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				13223 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				13227 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				13244 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				13250 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				13267 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				13271 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				13290 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				13350 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				13470 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				13517 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				13526 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				13532 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				13612 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				13634 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				13639 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				13666 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				13668 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				13714 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				13727 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				13756 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				13830 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				13838 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				13864 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				13938 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				13965 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				14010 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				14049 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				14092 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				14114 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				14186 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				14300 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				14339 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				14415 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				14419 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				14445 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				14453 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				14470 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				14501 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				14605 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				14667 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				14707 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				14720 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				14762 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				14781 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				14821 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				14850 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				14875 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				14904 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				14954 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				15048 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				15091 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				15093 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				15146 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				15163 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				15187 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				15206 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				15273 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				15393 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				15467 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				15481 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				15510 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				15625 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				15668 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				15679 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				15718 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				15769 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				15825 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				15860 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				15909 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				15947 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				15948 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				16125 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				16136 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				16194 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				16213 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				16354 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				16372 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				16480 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				16570 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				16586 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				16598 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				16725 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				16847 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				16862 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				16878 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				16912 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				16986 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				17003 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				17034 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				17092 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				17117 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				17147 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				17155 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				17166 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				17209 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				17233 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				17255 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				17360 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				17364 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				17387 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				17396 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				17404 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				17440 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				17466 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				17621 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				17691 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				17753 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				17774 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				17779 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				17806 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				17814 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				17846 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				17930 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				17951 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				17955 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				17966 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				17976 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				18001 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				18113 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				18257 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				18274 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				18283 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				18316 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				18324 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				18325 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				18372 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				18379 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				18395 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				18461 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				18475 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				18502 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				18504 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				18515 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				18561 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				18615 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				18618 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				18623 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				18681 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				18880 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				18953 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				18975 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				18999 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				19012 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				19021 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				19071 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				19072 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				19123 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				19157 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				19159 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				19171 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				19181 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				19314 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				19325 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				19329 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				19341 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				19414 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				19449 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				19461 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				19465 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				19469 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				19479 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				19539 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				19564 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				19609 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				19625 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				19633 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				19648 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				19653 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				19658 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				19700 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				19705 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				19713 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				19728 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				19729 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				19743 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				19761 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				19767 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				19795 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				19830 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				19915 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				19917 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				19951 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				19970 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				19972 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				19979 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				19995 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				19998 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				20016 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				20035 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				20105 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				20114 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				20124 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				20132 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				20202 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				20340 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				20348 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				20354 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				20382 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				20434 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				20441 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				20458 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				20472 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				20523 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				20527 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				20529 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				20537 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				20546 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				20587 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				20598 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				20627 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				20640 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				20686 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				20696 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				20713 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				20752 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				20760 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				20801 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				20861 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				20876 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				20927 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				20977 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				21011 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				21025 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				21052 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				21081 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				21092 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				21101 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				21215 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				21224 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				21244 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				21254 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				21268 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				21306 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				21310 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				21311 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				21356 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				21362 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				21371 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				21395 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				21406 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				21447 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				21470 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				21490 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				21523 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				21549 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				21587 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				21667 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				21678 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				21737 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				21880 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				21914 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				21951 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				21989 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				22004 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				22035 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				22036 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				22083 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				22152 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				22170 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				22177 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				22263 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				22299 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				22308 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				22333 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				22346 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				22356 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				22402 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				22412 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				22474 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				22483 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				22505 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				22512 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				22541 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				22602 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				22711 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				22765 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				22770 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				22779 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				22785 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				22815 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				22821 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				22852 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				22855 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				22934 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				22963 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				22970 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				22971 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				23025 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				23026 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				23054 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				23064 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				23067 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				23166 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				23233 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				23244 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				23259 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				23369 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				23416 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				23425 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				23497 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				23511 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				23512 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				23517 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				23558 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				23560 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				23586 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				23606 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				23609 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				23619 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				23620 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				23646 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				23647 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				23698 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				23706 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				23719 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				23771 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				23778 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				23793 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				23802 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				23816 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				23817 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				23861 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				23963 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				24063 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				24071 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				24079 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				24109 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				24120 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				24123 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				24155 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				24236 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				24264 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				24271 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				24305 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				24350 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				24352 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				24393 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				24404 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				24427 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				24436 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				24480 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				24484 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				24527 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				24546 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				24558 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				24559 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				24582 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				24654 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				24682 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				24774 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				24783 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				24807 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				24844 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				24931 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				24985 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				24991 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				25042 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				25047 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				25069 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				25108 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				25124 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				25160 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				25260 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				25383 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				25410 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				25427 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				25435 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				25500 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				25602 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				25651 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				25697 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				25698 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				25789 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				25824 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				25884 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				25898 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				25923 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				25952 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				25964 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				26053 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				26069 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				26131 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				26183 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				26229 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				26299 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				26319 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				26364 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				26376 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				26449 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				26583 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				26619 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				26649 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				26702 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				26772 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				26778 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				26784 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				26842 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				26846 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				26870 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				26895 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				26904 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				26941 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				26948 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				26988 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				27003 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				27033 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				27081 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				27087 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				27091 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				27290 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				27294 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				27377 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				27400 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				27451 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				27470 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				27486 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				27544 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				27579 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				27610 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				27625 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				27673 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				27731 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				27754 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				27767 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				27769 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				27781 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				27784 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				27800 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				27856 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				27903 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				27957 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				28014 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				28028 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				28034 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				28178 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				28192 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				28207 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				28259 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				28292 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				28296 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				28321 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				28402 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				28446 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				28471 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				28502 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				28552 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				28577 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				28627 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				28628 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				28652 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				28653 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				28682 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				28704 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				28716 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				28753 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				28758 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				28770 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				28783 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				28796 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				28826 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				28854 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				28861 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				28914 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				28915 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				28923 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				29027 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				29065 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				29070 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				29073 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				29097 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				29161 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				29177 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				29197 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				29229 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				29305 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				29330 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				29351 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				29375 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				29399 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				29418 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				29427 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				29438 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				29454 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				29511 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				29522 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				29561 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				29583 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				29609 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				29729 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				29812 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				29835 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				29887 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				30055 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				30083 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				30086 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				30135 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				30161 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				30162 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				30172 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				30194 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				30254 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				30316 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				30333 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				30347 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				30372 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				30385 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				30424 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				30487 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				30510 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				30557 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				30585 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				30664 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				30668 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				30681 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				30688 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				30720 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				30721 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				30739 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				30806 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				30862 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				30912 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				30945 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				30950 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				30953 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				30973 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				31001 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				31017 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				31083 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				31101 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				31176 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				31198 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				31213 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				31220 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				31222 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				31254 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				31256 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				31257 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				31315 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				31337 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				31353 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				31385 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				31392 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				31404 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				31499 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				31519 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				31529 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				31566 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				31617 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				31633 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				31700 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				31743 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				31884 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				31889 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				31904 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				31937 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				31953 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				32025 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				32042 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				32111 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				32212 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				32226 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				32247 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				32357 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				32371 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				32419 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				32420 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				32459 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				32495 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				32534 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				32581 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				32585 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				32637 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				32706 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				32715 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				32718 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				32732 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				32780 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				32793 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				32796 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				32809 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				32828 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				32885 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				32887 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				32959 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				32963 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				32968 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				32979 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				33090 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				33285 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				33337 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				33386 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				33408 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				33487 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				33571 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				33578 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				33608 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				33630 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				33637 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				33671 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				33677 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				33688 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				33747 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				33809 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				33810 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				33825 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				33834 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				33872 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				33914 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				33929 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				33949 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				33954 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				33971 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				33999 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				34029 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				34107 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				34122 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				34184 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				34231 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				34250 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				34298 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				34478 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				34606 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				34615 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				34623 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				34650 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				34673 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				34739 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				34798 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				34824 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				34888 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				34922 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				34924 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				35039 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				35045 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				35081 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				35120 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				35130 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				35140 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				35187 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				35207 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				35214 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				35240 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				35300 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				35305 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				35372 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				35373 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				35382 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				35388 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				35438 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				35447 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				35452 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				35485 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				35508 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				35510 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				35526 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				35575 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				35593 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				35596 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				35602 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				35670 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				35703 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				35748 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				35779 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				35784 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				35813 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				35864 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				35885 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				35888 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				35953 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				36012 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				36013 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				36024 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				36037 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				36073 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				36083 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				36108 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				36113 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				36141 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				36144 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				36156 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				36204 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				36282 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				36299 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				36313 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				36322 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				36351 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				36360 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				36435 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				36439 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				36467 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				36469 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				36506 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				36524 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				36559 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				36589 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				36638 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				36667 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				36706 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				36726 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				36751 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				36770 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				36801 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				36816 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				36841 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				36885 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				36933 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				36935 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				37105 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				37161 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				37162 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				37242 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				37244 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				37273 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				37364 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				37400 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				37421 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				37432 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				37508 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				37520 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				37528 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				37543 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				37562 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				37563 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				37682 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				37685 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				37714 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				37717 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				37718 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				37759 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				37766 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				37783 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				37872 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				37949 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				37961 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				38001 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				38054 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				38096 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				38138 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				38190 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				38297 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				38413 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				38461 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				38462 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				38503 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				38532 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				38563 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				38604 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				38631 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				38675 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				38681 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				38734 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				38761 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				38766 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				38791 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				38825 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				38836 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				38860 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				38911 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				38936 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				38962 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				39096 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				39117 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				39191 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				39200 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				39224 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				39267 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				39268 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				39297 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				39332 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				39377 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				39380 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				39425 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				39469 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				39482 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				39498 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				39590 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				39606 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				39621 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				39625 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				39719 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				39773 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				39779 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				39911 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				40042 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				40160 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				40162 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				40193 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				40261 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				40281 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				40343 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				40378 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				40457 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				40464 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				40532 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				40539 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				40543 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				40553 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				40559 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				40564 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				40632 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				40638 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				40645 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				40689 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				40713 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				40741 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				40803 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				40818 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				40885 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				40907 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				40943 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				40946 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				40951 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				40968 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				41024 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				41037 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				41076 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				41078 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				41121 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				41159 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				41200 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				41293 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				41320 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				41352 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				41372 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				41390 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				41424 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				41451 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				41509 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				41510 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				41555 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				41562 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				41670 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				41678 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				41701 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				41730 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				41816 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				41834 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				41848 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				41902 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				41903 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				41921 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				41934 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				41945 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				41946 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				42004 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				42016 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				42037 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				42040 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				42045 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				42089 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				42123 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				42161 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				42164 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				42213 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				42216 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				42344 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				42387 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				42456 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				42458 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				42554 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				42559 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				42562 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				42580 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				42636 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				42673 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				42719 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				42795 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				42847 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				42970 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				42992 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				42998 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				43065 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				43068 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				43072 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				43103 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				43140 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				43167 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				43180 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				43202 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				43306 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				43316 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				43385 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				43397 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				43401 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				43413 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				43439 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				43444 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				43470 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				43553 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				43557 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				43560 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				43581 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				43599 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				43622 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				43645 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				43667 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				43712 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				43782 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				43841 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				43843 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				43850 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				43856 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				43868 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				43869 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				43927 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				43930 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				43943 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				43953 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				43996 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				44044 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				44062 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				44121 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				44144 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				44166 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				44258 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				44390 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				44449 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				44606 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				44618 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				44619 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				44643 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				44673 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				44695 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				44765 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				44792 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				44810 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				44869 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				44914 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				44927 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				44947 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				44969 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				44994 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				45000 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				45051 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				45093 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				45114 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				45126 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				45135 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				45153 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				45165 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				45166 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				45168 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				45210 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				45266 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				45333 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				45401 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				45415 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				45440 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				45531 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				45549 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				45620 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				45665 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				45674 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				45780 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				45823 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				45848 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				45883 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				45909 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				45918 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				45933 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				45968 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				45972 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				45994 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				45998 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				46008 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				46048 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				46074 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				46079 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				46140 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				46164 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				46221 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				46237 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				46310 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				46312 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				46373 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				46468 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				46523 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				46528 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				46557 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				46576 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				46584 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				46599 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				46613 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				46661 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				46709 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				46789 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				46794 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				46803 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				46807 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				46810 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				46861 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				46867 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				46881 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				46887 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				46933 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				47007 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				47042 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				47078 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				47093 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				47106 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				47155 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				47176 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				47180 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				47183 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				47189 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				47223 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				47275 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				47279 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				47282 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				47290 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				47302 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				47344 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				47357 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				47398 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				47401 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				47579 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				47585 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				47602 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				47637 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				47647 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				47761 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				47915 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				47923 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				47935 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				47957 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				48031 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				48038 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				48062 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				48088 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				48097 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				48169 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				48173 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				48187 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				48192 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				48209 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				48211 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				48217 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				48219 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				48390 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				48404 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				48406 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				48414 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				48416 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				48433 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				48469 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				48480 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				48500 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				48529 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				48534 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				48541 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				48573 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				48638 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				48648 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				48650 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				48770 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				48775 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				48835 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				48870 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				48947 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				48967 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				48987 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				49098 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				49113 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				49120 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				49232 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				49241 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				49255 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				49322 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				49324 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				49443 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				49452 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				49479 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				49526 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				49539 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				49579 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				49610 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				49657 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				49671 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				49699 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				49734 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				49781 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				49802 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				49806 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				49870 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				49880 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				49911 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				49917 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				49948 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				49951 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				50031 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				50050 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				50054 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				50056 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				50145 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				50149 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				50274 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				50338 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				50386 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				50424 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				50434 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				50477 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				50495 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				50497 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				50504 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				50560 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				50659 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				50690 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				50711 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				50726 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				50772 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				50787 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				50860 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				50866 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				50921 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				50975 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				50983 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				51024 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				51036 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				51054 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				51059 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				51168 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				51206 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				51232 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				51244 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				51254 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				51328 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				51351 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				51363 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				51388 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				51400 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				51404 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				51436 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				51620 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				51633 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				51674 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				51759 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				51823 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				51837 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				51897 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				51958 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				52026 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				52157 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				52269 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				52278 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				52290 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				52392 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				52404 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				52418 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				52424 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				52439 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				52466 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				52481 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				52485 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				52495 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				52510 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				52523 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				52568 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				52570 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				52571 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				52575 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				52584 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				52776 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				52786 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				52882 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				52883 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				52893 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				52943 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				52947 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				52968 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				53002 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				53006 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				53023 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				53071 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				53074 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				53076 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				53101 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				53164 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				53167 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				53201 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				53220 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				53268 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				53292 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				53294 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				53317 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				53338 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				53399 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				53429 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				53460 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				53461 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				53500 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				53503 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				53523 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				53524 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				53539 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				53542 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				53565 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				53603 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				53641 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				53721 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				53732 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				53779 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				53830 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				53845 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				53922 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				53945 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				53958 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				53993 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				53998 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				54035 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				54054 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				54107 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				54118 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				54195 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				54196 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				54250 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				54254 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				54293 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				54300 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				54331 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				54416 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				54470 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				54494 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				54505 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				54526 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				54632 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				54714 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				54741 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				54780 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				54972 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				54977 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				54984 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				54987 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				54995 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				55012 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				55080 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				55109 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				55131 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				55165 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				55201 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				55277 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				55296 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				55301 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				55533 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				55608 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				55668 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				55785 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				55870 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				55914 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				55916 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				55937 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				56136 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				56176 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				56238 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				56239 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				56248 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				56258 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				56271 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				56343 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				56382 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				56384 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				56447 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				56508 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				56527 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				56547 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				56583 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				56703 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				56731 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				56783 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				56832 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				56835 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				56869 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				56897 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				56910 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				56927 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				56970 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				57030 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				57034 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				57074 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				57102 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				57107 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				57147 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				57167 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				57173 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				57179 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				57197 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				57203 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				57212 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				57251 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				57254 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				57304 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				57325 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				57341 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				57362 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				57373 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				57419 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				57448 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				57452 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				57475 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				57479 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				57490 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				57520 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				57530 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				57543 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				57593 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				57627 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				57632 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				57635 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				57749 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				57778 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				57835 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				57838 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				57844 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				57898 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				57943 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				57984 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				57991 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				58055 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				58215 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				58227 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				58263 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				58264 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				58300 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				58320 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				58346 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				58402 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				58531 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				58562 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				58606 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				58636 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				58699 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				58798 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				58889 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				58910 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				59054 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				59135 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				59156 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				59179 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				59182 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				59235 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				59330 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				59348 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				59372 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				59376 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				59596 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				59597 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				59628 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				59629 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				59695 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				59742 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				59745 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				59747 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				59767 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				59790 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				59792 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				59825 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				59826 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				59858 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				59901 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				59961 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				60032 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				60053 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				60058 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				60068 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				60071 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				60128 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				60130 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				60184 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				60250 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				60264 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				60298 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				60299 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				60497 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				60498 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				60550 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				60618 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				60679 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				60688 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				60691 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				60791 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				60903 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				60917 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				60929 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				60930 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				60951 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				60963 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				60964 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				60967 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				61061 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				61130 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				61133 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				61159 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				61185 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				61220 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				61227 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				61267 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				61293 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				61313 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				61388 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				61425 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				61488 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				61542 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				61595 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				61596 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				61635 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				61769 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				61775 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				61805 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				61816 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				62033 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				62070 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				62081 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				62190 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				62299 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				62321 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				62328 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				62361 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				62382 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				62389 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				62454 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				62469 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				62491 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				62531 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				62534 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				62542 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				62610 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				62645 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				62655 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				62668 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				62711 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				62740 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				62802 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				62823 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				62845 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				62851 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				62935 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				62993 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				63053 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				63099 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				63101 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				63109 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				63221 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				63287 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				63289 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				63291 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				63311 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				63327 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				63374 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				63409 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				63691 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				63712 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				63775 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				63785 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				63811 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				63822 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				63842 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				63854 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				63884 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				63903 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				63914 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				63933 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				63976 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				64005 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				64014 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				64049 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				64111 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				64118 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				64144 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				64158 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				64189 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				64195 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				64289 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				64361 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				64372 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				64407 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				64442 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				64458 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				64491 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				64496 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				64514 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				64516 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				64636 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				64659 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				64713 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				64727 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				64751 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				64782 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				64814 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				64816 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				64824 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				64825 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				64839 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				64844 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				64855 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				64876 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				64903 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				64960 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				65011 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				65043 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				65147 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				65178 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				65186 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				65278 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				65306 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				65338 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				65367 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				65369 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				65375 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				65477 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				65478 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),

                                OTHERS => STD_LOGIC_VECTOR(to_unsigned(238, 8))
                            );
                    
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
                ASSERT (mem_we = '1' OR mem_we = '0') REPORT "o_mem_we in an unexpected state" SEVERITY failure;
            END IF;
            ASSERT (enable_wire = '1' OR enable_wire = '0') REPORT "o_mem_en in an unexpected state" SEVERITY failure;
        END IF;
    END PROCESS;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    createScenario : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '0' THEN
            tb_rst <= scenario_rst(0);
            tb_w <= scenario_w(0);
            tb_start <= scenario_start(0);
            scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_done = '0' REPORT "TEST FALLITO (postreset DONE != 0 )" SEVERITY failure;
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0001110011100111:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0011000100010111:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0010100111011011:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(133, 8)) severity failure; -- 1111110100101111:133->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 000111000000001:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 01111100100011:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0001111001000001:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1100101110001:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1000101011011:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1011101100011:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 001000110101101:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(243, 8)) severity failure; -- 0100010101111111:243->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(243, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0001001001010101:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(243, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1001101000110011:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0101100101000101:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 11111001000011:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 11110010011:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0100000000000111:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0011001110110101:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1010101001001111:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0010110101010101:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1000001110101111:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0011000000111111:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 001111100111001:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 10000001011101:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1101011110011101:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 110100000111111:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1000100111100101:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0110111110011111:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 01001110100111:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0100111110110111:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0101000100111:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0101100111111011:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 001110110101001:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0111110101110011:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 101100110110101:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 10001000001111:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 000110101010011:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0111100111010001:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0111101011001:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0000101001111001:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0001100111101111:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 110011000100111:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1100010001001011:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 10011001100011:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0011110010110111:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1000011111010101:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 00001100110011:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 010100000000101:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0010010010100111:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 001110101110111:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 000000010001101:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0011110001011101:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 100101001001011:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1110001101001111:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 11100010111101:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 101001011000001:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1001001011101101:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0000010100100111:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1001001100101111:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 11011000000101:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1100001001100001:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0111100000111:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0101010010101011:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 10000000001:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 00000000000011:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 001000011001001:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0110110010100111:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0001000001101011:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0010100000010111:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 111100010110101:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 010100100100001:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 11011101011111:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1111000111000011:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0111100101110101:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 10010010110001:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1001001001101011:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0110011101111:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 111011101100101:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 011100111011101:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1101010100100011:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1000001001110101:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 00000101010001:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8)) severity failure; -- 0011111000111111:108->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 000011111110011:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1000101101101001:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 001100000011:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 01101011110011:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1011110001111111:238->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1010100011110111:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 1101010010001011:238->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 101000010111:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 0011000100101:238->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- 111101010001001:238->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 

        ASSERT false REPORT "Simulation Ended! TEST PASSATO (EXAMPLE)" SEVERITY failure;
    END PROCESS testRoutine;

END projecttb;
