LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 2801; 
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00110" & "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000" & "111111111111111111000011111111111111111100000000000000011111111111111111000000000000000000000000000000011111111111111111000000011111111111111111100000000000000000011111111111111111100000000001111111111111111100000000000000000000000000000001111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111110000000011111111111111111100000000000000000000000000000011111111111111111100000000000000000000000000000111111111111111100000000000000000000000000000011111111111111111000000000000000000000000000000111111111111111111000000000000000000000000001111111111111111000000000000011111111111111110000000000111111111111111111000000000000000000000000000001111111111111111110000000011111111111111111100000000000000000000111111111111111111000000000000000000000000000000111111111111111111000000000000111111111111111111000000000000000000000011111111111111111000000000000111111111111111111000000000000000000000000001111111111111111100000000000000000011111111111111111100000000000000000111111111111111111000000000000000111111111111111111000000000000000000000000111111111111110000000000000000000000000000000111111111111111111000000000000000000111111111111111000000000000000000000000001111111111111111100000111111111111111111000000000000000000000000000000111111111111111111000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000000011111111111111111100000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000000000111111111111111111000000000000000000000011111111111111111100000011111111111111111000001111111111111111100000000000111111111111111111000000000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000001111111111111111110000000000111111111111111111000000000000000000000000000011111111111111111000000000000111111111111111111000000111111111111111110000000000000011111111111111111100000000000011111111111111111100000000000000000111111111111111111000000000000000000000000000011111111111111111100000000000000000000000000001111111111111111110000000000000001111111111111111110000000111111111111111000000000000000000000001111111111111111110000000111111111111111111000000000000011111111111111111100000000000000001111111111111111110000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000011111111111111100000000000011111111111111111100000011111111111111111100000000000000000111111111111110000000000000000000000001111111111111111110000000000000000000000000000000111111111111111111000000000000000";
    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000" & "000110011101110111000000011000010001000100000000000000010001000111110111000000000000000000000000000000001000111110001111000000011111001010011100100000000000000000010101001001110100100000000001101101111101111100000000000000000000000000000001111000010010000000000000000000000110110010010100011000000000000000000000000011101101110000110000000011101000110111100100000000000000000000000000000000101001111010010100000000000000000000000000000010001000101000100000000000000000000000000000011010101100100001000000000000000000000000000000001000010110001111000000000000000000000000001110000101111001000000000000001111010111011110000000000110001101110000001000000000000000000000000000000111111001001000110000000010000001111001101100000000000000000000110010111000001101000000000000000000000000000000111001001001110111000000000000001010001110110111000000000000000000000011101111001110011000000000000110111010101101101000000000000000000000000001111110000010011100000000000000000011011100011010011100000000000000000111110001011010111000000000000000001101001001100001000000000000000000000000011001111101010000000000000000000000000000000111110101010101111000000000000000000111011000001011000000000000000000000000000100001010000010100000100101101010110001000000000000000000000000000000011110111111111101000000000000111111100011001011000000000000000000000000001000010111100010100000000000000000000000000011000001111100000100000000011100111010011011000000000000000000000000110101010101010001000000000000000000000000000000101100010001110101000000000000000000000001101010011001001100000010001101010011011000000011011100001100100000000000111111010000101111000000000000000000000000000000101101111001001001000000000000000000000000010001011001011100000000000000000010001011011111000100000000000000000000000001000011100111010000000000000000001100100001000010110000000000100010010111110111000000000000000000000000000011111011011100001000000000000111001000111010001000000111011101100100010000000000000000110111010111100100000000000001000110011011000100000000000000000110000110001000101000000000000000000000000000010000000010011010100000000000000000000000000000000100111010000110000000000000001100111011000001010000000000100110101001000000000000000000000001001000001011010010000000111001101101111001000000000000011010011111011100100000000000000000001111110100000010000000000000000110110101110101001000000000000000000000011111000000101011100000000000000000000000000001001101010100111100000000000000000000000011000010010111011100000000000000000000000001111011101100011100000000000000000000001000010101100010000000000000000011100101010101100000000000011111011100000100100000001010101110000111100000000000000000111001100111010000000000000000000000000110110001011100110000000000000000000000000000000011100000101111011000000000000000";

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (  
				23 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				144 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				162 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				179 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				194 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				282 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				329 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				330 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				339 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				362 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				445 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				482 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				484 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				490 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				564 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				684 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				691 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				708 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				713 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				730 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				752 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				809 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				823 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				872 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				902 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				904 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				937 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				943 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				985 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				997 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				1016 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				1023 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				1037 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				1143 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				1152 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				1176 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				1302 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				1308 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				1368 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				1384 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				1389 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				1458 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				1459 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				1505 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				1534 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				1575 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				1594 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				1625 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				1646 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				1647 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				1710 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				1730 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				1807 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				1848 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				1862 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				1899 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				1945 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				1949 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				1960 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				1963 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				1989 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				2024 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				2027 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				2029 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				2108 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				2122 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				2143 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				2150 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				2174 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				2240 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				2250 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				2291 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				2365 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				2446 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				2493 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				2546 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				2575 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				2611 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				2651 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				2713 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				2740 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				2742 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				2768 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				2894 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				2915 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				2928 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				2942 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				2949 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				2975 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				3009 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				3061 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				3098 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				3099 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				3120 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				3134 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				3176 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				3190 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				3225 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				3235 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				3272 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				3335 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				3365 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				3367 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				3448 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				3500 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				3522 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				3582 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				3586 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				3694 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				3725 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				3728 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				3756 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				3777 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				3797 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				3823 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				3828 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				3841 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				3963 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				3964 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				3972 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				4001 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				4004 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				4024 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				4036 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				4093 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				4126 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				4171 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				4218 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				4244 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				4299 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				4362 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				4366 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				4387 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				4389 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				4411 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				4535 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				4560 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				4599 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				4631 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				4640 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				4660 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				4681 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				4687 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				4690 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				4702 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				4715 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				4785 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				4824 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				4853 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				4895 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				4977 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				4993 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				4995 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				5039 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				5042 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				5048 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				5156 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				5178 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				5196 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				5240 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				5358 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				5387 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				5436 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				5467 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				5484 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				5680 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				5804 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				5841 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				5842 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				5967 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				6033 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				6130 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				6166 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				6192 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				6212 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				6213 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				6282 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				6296 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				6359 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				6432 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				6461 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				6472 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				6534 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				6547 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				6556 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				6598 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				6600 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				6711 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				6736 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				6754 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				6902 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				6926 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				6961 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				6999 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				7025 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				7032 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				7054 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				7071 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				7110 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				7176 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				7205 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				7236 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				7273 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				7293 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				7298 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				7304 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				7332 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				7339 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				7374 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				7378 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				7412 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				7422 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				7495 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				7551 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				7619 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				7737 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				7775 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				7786 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				7874 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				7896 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				8081 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				8094 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				8131 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				8165 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				8222 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				8234 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				8236 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				8254 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				8257 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				8294 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				8312 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				8330 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				8391 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				8402 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				8421 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				8447 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				8449 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				8502 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				8544 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				8570 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				8573 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				8611 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				8614 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				8615 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				8642 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				8647 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				8648 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				8679 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				8762 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				8777 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				8808 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				8820 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				8822 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				8883 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				8963 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				8965 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				8994 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				9022 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				9140 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				9156 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				9166 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				9186 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				9190 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				9198 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				9203 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				9215 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				9255 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				9259 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				9275 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				9301 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				9322 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				9345 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				9398 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				9491 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				9500 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				9589 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				9652 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				9670 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				9687 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				9738 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				9786 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				9799 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				9825 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				9968 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				10005 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				10035 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				10046 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				10102 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				10153 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				10162 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				10200 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				10206 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				10222 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				10248 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				10287 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				10294 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				10390 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				10431 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				10451 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				10477 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				10491 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				10565 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				10642 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				10656 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				10691 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				10711 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				10849 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				10864 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				10877 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				10952 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				10959 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				10970 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				11003 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				11049 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				11102 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				11205 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				11225 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				11233 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				11261 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				11268 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				11282 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				11292 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				11303 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				11338 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				11416 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				11483 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				11502 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				11563 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				11617 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				11664 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				11669 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				11698 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				11836 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				11850 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				11863 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				11988 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				12036 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				12045 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				12069 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				12071 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				12080 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				12102 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				12154 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				12208 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				12266 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				12276 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				12297 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				12318 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				12326 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				12328 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				12460 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				12487 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				12598 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				12599 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				12624 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				12660 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				12670 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				12679 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				12773 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				12797 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				12840 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				12850 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				12951 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				12978 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				13018 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				13031 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				13116 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				13132 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				13133 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				13134 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				13177 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				13199 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				13233 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				13267 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				13314 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				13317 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				13329 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				13344 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				13356 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				13456 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				13489 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				13491 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				13514 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				13635 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				13708 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				13817 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				13861 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				13882 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				13887 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				13891 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				13938 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				14019 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				14042 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				14044 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				14096 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				14164 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				14199 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				14206 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				14212 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				14219 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				14245 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				14258 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				14276 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				14390 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				14399 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				14401 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				14410 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				14414 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				14425 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				14427 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				14437 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				14518 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				14575 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				14628 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				14669 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				14720 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				14729 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				14774 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				14824 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				14850 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				14889 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				14902 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				14926 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				14945 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				15126 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				15181 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				15222 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				15250 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				15264 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				15265 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				15266 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				15334 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				15413 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				15468 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				15484 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				15533 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				15545 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				15567 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				15568 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				15597 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				15709 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				15738 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				15766 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				15829 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				15833 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				15854 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				15878 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				15929 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				15934 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				15947 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				15980 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				15984 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				15988 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				16015 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				16085 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				16099 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				16120 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				16179 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				16313 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				16349 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				16390 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				16407 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				16452 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				16499 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				16619 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				16654 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				16658 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				16737 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				16742 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				16786 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				16811 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				16922 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				16946 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				17021 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				17030 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				17040 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				17056 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				17077 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				17118 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				17137 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				17156 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				17227 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				17248 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				17267 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				17311 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				17331 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				17360 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				17391 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				17396 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				17425 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				17492 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				17523 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				17527 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				17589 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				17631 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				17632 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				17698 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				17805 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				17841 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				17884 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				17901 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				17903 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				17921 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				17953 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				17986 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				18004 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				18041 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				18119 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				18123 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				18134 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				18150 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				18157 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				18183 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				18221 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				18431 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				18485 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				18506 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				18517 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				18610 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				18615 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				18659 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				18676 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				18714 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				18726 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				18757 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				18771 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				18776 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				18851 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				18858 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				18990 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				18994 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				19036 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				19040 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				19090 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				19093 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				19106 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				19125 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				19149 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				19165 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				19187 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				19244 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				19344 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				19359 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				19388 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				19401 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				19423 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				19437 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				19590 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				19605 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				19780 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				19851 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				19879 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				20127 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				20128 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				20129 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				20355 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				20477 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				20493 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				20519 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				20573 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				20598 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				20623 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				20648 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				20650 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				20663 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				20686 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				20734 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				20751 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				20773 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				20816 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				20892 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				20902 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				20983 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				21042 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				21078 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				21351 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				21360 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				21391 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				21413 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				21471 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				21521 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				21532 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				21535 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				21544 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				21560 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				21595 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				21635 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				21657 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				21662 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				21664 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				21674 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				21689 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				21789 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				21842 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				21850 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				21851 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				21867 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				21944 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				21994 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				21997 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				22043 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				22064 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				22084 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				22139 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				22166 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				22231 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				22271 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				22306 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				22431 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				22436 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				22440 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				22442 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				22575 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				22605 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				22657 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				22695 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				22698 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				22703 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				22715 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				22721 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				22788 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				22821 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				22839 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				22844 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				22852 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				22898 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				22923 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				22982 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				23034 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				23063 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				23115 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				23124 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				23125 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				23161 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				23168 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				23199 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				23219 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				23242 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				23282 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				23392 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				23422 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				23442 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				23470 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				23476 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				23529 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				23562 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				23566 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				23614 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				23667 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				23682 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				23757 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				23787 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				23827 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				23852 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				23899 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				23907 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				23934 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				23938 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				23942 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				24052 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				24126 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				24156 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				24166 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				24299 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				24349 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				24355 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				24391 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				24408 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				24438 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				24442 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				24447 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				24448 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				24455 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				24501 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				24502 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				24525 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				24574 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				24649 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				24673 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				24676 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				24684 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				24704 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				24789 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				24827 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				24864 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				24893 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				24896 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				24994 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				25017 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				25251 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				25290 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				25363 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				25400 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				25425 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				25434 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				25452 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				25485 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				25644 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				25647 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				25700 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				25701 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				25730 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				25774 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				25781 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				25790 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				25803 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				25833 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				25873 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				25893 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				25942 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				25992 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				26023 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				26033 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				26048 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				26067 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				26069 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				26080 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				26107 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				26146 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				26185 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				26188 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				26211 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				26287 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				26311 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				26329 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				26365 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				26421 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				26505 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				26512 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				26529 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				26546 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				26603 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				26652 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				26659 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				26665 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				26705 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				26729 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				26745 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				26789 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				26792 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				26793 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				26804 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				26978 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				26989 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				26995 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				27024 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				27062 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				27100 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				27117 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				27124 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				27143 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				27299 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				27386 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				27426 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				27453 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				27497 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				27579 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				27583 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				27609 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				27702 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				27708 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				27714 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				27731 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				27745 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				27869 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				27880 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				27885 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				27926 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				27927 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				27968 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				28018 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				28151 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				28227 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				28268 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				28390 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				28406 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				28410 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				28502 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				28535 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				28550 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				28584 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				28595 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				28643 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				28766 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				28770 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				28867 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				28868 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				28904 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				28921 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				28928 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				28950 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				28974 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				28992 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				28996 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				29052 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				29063 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				29086 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				29136 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				29179 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				29186 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				29229 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				29241 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				29309 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				29333 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				29334 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				29404 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				29459 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				29472 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				29502 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				29527 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				29536 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				29578 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				29579 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				29625 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				29669 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				29710 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				29760 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				29793 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				29797 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				29798 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				29824 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				29830 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				29855 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				29886 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				29917 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				29921 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				29992 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				30015 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				30050 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				30074 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				30252 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				30283 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				30292 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				30379 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				30442 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				30581 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				30592 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				30593 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				30843 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				30901 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				30931 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				30941 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				30956 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				30964 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				31000 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				31051 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				31080 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				31111 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				31152 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				31155 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				31244 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				31304 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				31322 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				31394 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				31722 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				31740 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				31743 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				31783 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				31860 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				31879 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				31920 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				31929 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				31931 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				31937 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				31949 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				32018 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				32084 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				32183 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				32190 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				32310 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				32425 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				32461 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				32482 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				32573 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				32597 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				32610 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				32630 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				32697 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				32764 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				32770 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				32771 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				32800 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				32843 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				32846 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				32908 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				32946 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				32954 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				32975 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				32997 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				33003 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				33005 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				33056 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				33122 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				33131 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				33132 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				33201 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				33235 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				33355 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				33358 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				33400 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				33438 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				33452 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				33480 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				33520 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				33570 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				33586 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				33611 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				33726 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				33779 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				33797 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				33825 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				33840 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				33849 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				33886 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				33940 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				34013 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				34032 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				34106 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				34108 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				34161 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				34183 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				34284 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				34293 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				34312 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				34332 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				34353 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				34390 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				34431 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				34438 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				34492 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				34494 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				34521 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				34566 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				34592 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				34598 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				34609 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				34703 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				34727 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				34759 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				34812 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				34848 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				34916 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				34966 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				34982 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				35009 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				35092 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				35099 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				35111 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				35225 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				35316 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				35329 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				35370 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				35416 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				35434 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				35508 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				35609 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				35631 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				35634 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				35692 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				35720 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				35813 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				35863 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				35880 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				35918 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				35933 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				36106 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				36110 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				36148 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				36244 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				36301 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				36303 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				36312 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				36330 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				36377 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				36456 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				36487 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				36520 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				36528 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				36535 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				36559 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				36656 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				36673 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				36695 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				36762 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				36789 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				36803 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				36834 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				36860 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				36875 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				37009 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				37179 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				37261 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				37343 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				37346 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				37382 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				37414 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				37511 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				37563 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				37566 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				37599 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				37618 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				37625 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				37671 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				37683 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				37717 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				37723 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				37725 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				37757 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				37761 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				37787 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				37794 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				37803 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				37870 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				37892 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				37908 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				37956 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				37969 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				37979 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				38025 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				38066 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				38140 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				38196 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				38328 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				38376 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				38412 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				38439 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				38447 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				38473 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				38642 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				38656 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				38669 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				38704 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				38712 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				38721 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				38769 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				38828 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				38866 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				38876 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				38914 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				38930 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				38944 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				38953 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				38967 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				38992 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				39033 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				39036 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				39074 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				39080 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				39099 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				39149 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				39177 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				39215 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				39295 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				39345 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				39349 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				39430 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				39454 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				39462 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				39485 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				39489 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				39590 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				39667 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				39689 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				39785 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				39807 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				39833 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				39844 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				39903 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				39910 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				39952 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				39969 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				40008 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				40042 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				40058 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				40095 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				40173 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				40174 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				40196 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				40256 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				40283 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				40327 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				40330 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				40400 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				40555 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				40620 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				40645 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				40669 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				40696 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				40798 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				40818 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				40863 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				40914 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				40987 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				41015 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				41017 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				41018 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				41029 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				41032 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				41100 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				41103 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				41105 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				41123 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				41189 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				41193 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				41201 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				41212 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				41214 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				41284 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				41298 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				41305 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				41321 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				41334 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				41392 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				41395 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				41396 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				41412 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				41437 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				41505 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				41515 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				41521 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				41533 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				41543 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				41556 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				41600 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				41741 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				41761 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				41789 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				41832 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				41838 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				41881 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				41950 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				41959 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				41966 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				41977 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				41985 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				42158 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				42214 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				42249 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				42262 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				42270 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				42394 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				42413 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				42474 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				42569 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				42575 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				42604 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				42633 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				42679 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				42791 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				42946 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				43008 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				43107 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				43139 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				43242 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				43285 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				43291 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				43292 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				43329 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				43375 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				43428 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				43437 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				43563 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				43607 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				43689 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				43733 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				43806 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				43813 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				43814 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				43818 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				43835 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				43837 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				43870 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				43890 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				43900 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				44004 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				44008 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				44020 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				44030 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				44056 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				44060 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				44119 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				44139 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				44211 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				44283 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				44287 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				44293 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				44303 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				44307 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				44359 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				44393 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				44417 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				44425 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				44450 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				44498 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				44513 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				44606 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				44758 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				44769 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				44866 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				44885 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				44934 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				44948 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				45023 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				45034 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				45089 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				45097 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				45105 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				45135 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				45144 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				45148 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				45182 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				45185 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				45186 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				45198 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				45217 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				45218 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				45301 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				45332 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				45346 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				45591 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				45651 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				45691 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				45728 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				45802 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				45839 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				45846 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				45983 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				46005 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				46096 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				46128 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				46166 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				46183 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				46221 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				46248 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				46308 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				46311 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				46364 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				46375 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				46402 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				46407 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				46427 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				46488 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				46526 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				46548 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				46592 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				46627 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				46633 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				46638 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				46663 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				46680 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				46697 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				46773 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				46827 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				46843 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				46864 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				46910 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				46924 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				46970 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				47006 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				47019 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				47040 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				47174 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				47177 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				47213 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				47222 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				47325 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				47330 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				47394 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				47421 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				47433 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				47437 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				47455 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				47471 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				47476 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				47495 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				47598 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				47668 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				47718 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				47724 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				47743 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				47779 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				47831 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				47956 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				47984 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				48010 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				48017 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				48039 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				48062 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				48136 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				48204 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				48225 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				48245 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				48256 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				48279 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				48289 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				48303 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				48322 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				48328 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				48422 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				48431 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				48478 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				48546 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				48565 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				48684 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				48854 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				48909 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				48946 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				48957 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				48983 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				49000 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				49001 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				49035 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				49170 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				49171 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				49177 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				49273 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				49276 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				49306 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				49349 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				49358 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				49359 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				49445 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				49457 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				49517 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				49533 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				49661 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				49679 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				49690 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				49747 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				49801 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				49890 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				49956 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				50039 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				50174 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				50187 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				50196 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				50202 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				50238 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				50241 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				50284 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				50367 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				50394 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				50400 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				50416 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				50455 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				50507 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				50565 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				50585 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				50648 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				50654 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				50725 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				50794 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				50821 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				50822 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				50840 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				50906 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				50928 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				50939 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				51004 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				51031 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				51056 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				51083 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				51155 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				51174 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				51188 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				51209 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				51211 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				51276 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				51305 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				51360 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				51420 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				51461 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				51519 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				51618 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				51707 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				51758 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				51759 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				51774 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				51792 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				51826 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				51857 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				51949 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				52010 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				52080 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				52117 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				52153 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				52210 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				52218 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				52219 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				52224 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				52412 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				52463 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				52499 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				52502 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				52593 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				52629 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				52667 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				52724 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				52745 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				52752 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				52757 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				52816 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				52854 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				52921 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				52933 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				53011 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				53038 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				53039 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				53071 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				53247 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				53276 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				53356 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				53427 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				53574 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				53608 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				53647 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				53668 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				53799 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				53835 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				53941 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				54003 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				54013 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				54058 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				54062 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				54089 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				54101 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				54130 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				54190 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				54201 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				54208 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				54259 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				54296 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				54319 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				54404 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				54425 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				54445 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				54451 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				54478 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				54481 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				54504 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				54525 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				54529 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				54609 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				54664 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				54741 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				54746 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				54770 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				54813 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				54917 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				54963 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				54969 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				54978 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				55115 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				55140 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				55158 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				55193 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				55197 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				55222 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				55248 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				55284 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				55363 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				55424 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				55438 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				55494 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				55506 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				55532 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				55535 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				55885 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				55893 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				55947 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				55969 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				55992 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				56071 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				56161 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				56221 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				56325 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				56411 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				56435 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				56493 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				56562 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				56565 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				56568 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				56593 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				56726 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				56816 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				56886 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				56898 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				56918 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				56919 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				57071 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				57135 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				57295 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				57306 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				57318 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				57333 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				57361 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				57372 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				57383 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				57400 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				57435 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				57436 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				57443 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				57450 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				57519 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				57614 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				57616 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				57698 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				57732 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				57852 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				57882 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				57917 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				57988 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				57990 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				57997 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				58052 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				58110 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				58121 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				58137 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				58152 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				58172 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				58216 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				58243 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				58398 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				58410 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				58419 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				58481 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				58493 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				58666 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				58668 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				58700 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				58731 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				58805 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				58858 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				58895 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				59012 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				59019 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				59024 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				59026 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				59087 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				59095 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				59117 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				59223 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				59225 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				59239 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				59242 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				59276 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				59280 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				59327 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				59356 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				59390 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				59423 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				59497 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				59504 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				59512 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				59514 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				59551 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				59602 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				59603 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				59620 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				59625 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				59653 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				59700 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				59718 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				59731 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				59767 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				59810 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				59855 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				59888 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				59949 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				59955 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				60100 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				60132 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				60184 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				60203 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				60215 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				60237 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				60246 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				60259 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				60271 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				60293 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				60314 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				60331 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				60360 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				60516 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				60524 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				60533 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				60596 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				60684 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				60714 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				60747 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				60751 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				60809 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				60832 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				60853 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				60887 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				60896 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				60913 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				60961 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				61010 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				61047 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				61105 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				61108 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				61155 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				61276 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				61301 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				61384 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				61449 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				61528 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				61548 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				61573 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				61577 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				61605 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				61629 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				61717 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				61723 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				61745 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				61762 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				61763 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				61767 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				61850 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				61865 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				61922 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				61947 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				61987 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				62009 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				62032 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				62108 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				62148 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				62164 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				62201 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				62216 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				62217 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				62257 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				62314 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				62496 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				62557 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				62709 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				62754 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				62786 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				62844 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				62882 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				62884 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				62896 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				62966 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				63027 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				63116 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				63125 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				63131 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				63180 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				63210 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				63227 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				63248 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				63259 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				63294 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				63342 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				63387 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				63395 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				63401 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				63408 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				63437 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				63454 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				63459 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				63501 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				63534 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				63595 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				63626 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				63666 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				63676 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				63677 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				63678 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				63691 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				63706 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				63713 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				63721 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				63734 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				63787 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				63837 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				63955 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				63958 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				63985 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				64018 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				64034 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				64090 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				64135 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				64172 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				64244 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				64257 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				64263 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				64287 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				64325 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				64342 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				64411 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				64419 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				64464 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				64521 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				64542 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				64546 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				64577 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				64598 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				64642 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				64723 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				64737 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				64860 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				64909 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				64967 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				64978 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				64997 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				64998 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				65083 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				65164 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				65194 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				65234 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				65261 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				65282 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				65354 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),

                                OTHERS => STD_LOGIC_VECTOR(to_unsigned(125, 8)
                            );
                    
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
                ASSERT (mem_we = '1' OR mem_we = '0') REPORT "o_mem_we in an unexpected state" SEVERITY failure;
            END IF;
            ASSERT (enable_wire = '1' OR enable_wire = '0') REPORT "o_mem_en in an unexpected state" SEVERITY failure;
        END IF;
    END PROCESS;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    createScenario : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '0' THEN
            tb_rst <= scenario_rst(0);
            tb_w <= scenario_w(0);
            tb_start <= scenario_start(0);
            scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_done = '0' REPORT "TEST FALLITO (postreset DONE != 0 )" SEVERITY failure;
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8)) severity failure;	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 

        ASSERT false REPORT "Simulation Ended! TEST PASSATO (EXAMPLE)" SEVERITY failure;
    END PROCESS testRoutine;

END projecttb;