LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 188; 
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00110" & "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000" & "111111111111111111011111111111111111100111111111111100111111111111111110001111111111111111110001111111111111111000111111111111100111111111111111111111111111111110000111111111111111110";
    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000" & "100001100111011101001100101001110110100101010101100100010101011110100010000011010001010010010000110100101111011000011110111100100001010010110010100101100011110110000010001100111000110";

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (  
				19 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				52 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				59 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				74 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				79 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				100 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				188 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				203 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				272 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				278 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				292 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				294 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				325 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				365 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				399 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				401 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				437 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				547 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				696 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				697 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				719 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				749 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				794 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				880 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				912 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				959 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				969 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				1002 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				1042 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				1095 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				1101 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				1109 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				1133 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				1142 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				1159 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				1171 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				1231 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				1246 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				1413 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				1421 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				1422 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				1429 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				1434 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				1438 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				1504 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				1518 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				1618 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				1694 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				1884 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				1908 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				2060 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				2074 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				2124 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				2126 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				2129 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				2157 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				2160 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				2164 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				2204 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				2206 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				2250 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				2287 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				2355 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				2370 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				2380 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				2425 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				2441 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				2463 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				2464 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				2495 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				2496 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				2501 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				2528 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				2538 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				2543 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				2601 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				2672 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				2698 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				2740 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				2750 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				2850 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				2867 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				2950 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				2952 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				3013 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				3027 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				3049 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				3091 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				3097 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				3168 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				3169 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				3171 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				3216 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				3227 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				3229 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				3265 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				3285 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				3353 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				3372 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				3374 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				3377 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				3506 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				3525 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				3591 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				3607 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				3655 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				3661 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				3698 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				3735 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				3784 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				3834 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				3910 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				3917 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				3944 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				3958 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				3977 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				4004 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				4031 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				4053 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				4199 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				4208 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				4252 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				4256 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				4271 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				4319 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				4327 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				4329 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				4396 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				4467 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				4583 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				4655 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				4669 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				4699 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				4716 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				4873 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				4897 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				4931 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				4969 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				4978 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				4989 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				5007 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				5050 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				5052 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				5075 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				5082 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				5097 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				5136 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				5165 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				5321 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				5352 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				5380 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				5383 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				5387 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				5388 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				5450 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				5524 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				5556 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				5575 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				5609 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				5633 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				5649 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				5680 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				5681 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				5692 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				5703 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				5785 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				5787 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				5900 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				6005 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				6018 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				6030 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				6036 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				6089 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				6118 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				6121 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				6231 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				6285 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				6307 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				6364 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				6368 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				6380 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				6413 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				6437 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				6465 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				6503 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				6643 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				6651 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				6690 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				6698 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				6743 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				6752 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				6753 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				6778 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				6851 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				6905 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				6947 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				6956 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				6979 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				7005 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				7055 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				7064 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				7077 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				7115 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				7120 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				7128 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				7154 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				7237 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				7257 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				7362 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				7371 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				7396 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				7436 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				7451 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				7463 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				7503 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				7515 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				7520 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				7525 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				7563 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				7605 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				7673 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				7782 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				7806 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				8015 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				8034 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				8049 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				8050 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				8129 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				8132 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				8142 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				8182 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				8267 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				8332 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				8338 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				8350 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				8355 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				8418 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				8422 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				8476 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				8504 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				8537 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				8558 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				8561 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				8563 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				8691 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				8770 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				8783 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				8806 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				8853 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				8919 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				8991 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				9030 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				9111 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				9142 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				9147 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				9161 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				9264 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				9294 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				9307 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				9323 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				9341 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				9387 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				9451 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				9467 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				9509 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				9548 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				9566 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				9596 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				9622 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				9661 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				9662 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				9663 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				9698 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				9704 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				9774 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				9778 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				9786 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				9817 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				9855 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				9884 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				9960 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				9988 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				10008 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				10034 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				10048 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				10056 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				10066 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				10147 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				10205 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				10221 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				10268 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				10392 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				10444 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				10459 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				10500 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				10596 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				10637 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				10655 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				10695 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				10700 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				10728 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				10743 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				10751 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				10783 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				10802 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				10848 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				10859 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				10940 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				11042 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				11119 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				11210 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				11230 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				11245 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				11279 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				11336 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				11348 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				11383 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				11413 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				11427 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				11478 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				11488 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				11507 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				11528 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				11538 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				11554 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				11559 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				11564 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				11614 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				11625 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				11795 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				11799 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				11817 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				11883 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				11887 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				11978 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				12001 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				12016 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				12113 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				12158 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				12171 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				12202 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				12368 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				12370 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				12377 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				12451 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				12541 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				12566 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				12620 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				12623 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				12634 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				12662 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				12667 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				12695 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				12700 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				12705 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				12727 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				12737 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				12752 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				12773 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				12816 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				12837 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				12916 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				12937 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				12949 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				13073 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				13079 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				13081 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				13090 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				13133 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				13151 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				13157 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				13170 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				13208 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				13227 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				13258 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				13280 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				13341 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				13353 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				13372 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				13551 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				13597 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				13601 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				13619 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				13620 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				13631 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				13685 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				13764 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				13780 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				13781 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				13830 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				13952 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				13974 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				13990 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				13991 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				14093 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				14100 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				14120 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				14134 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				14136 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				14147 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				14150 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				14203 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				14214 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				14243 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				14281 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				14293 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				14361 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				14419 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				14421 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				14520 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				14552 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				14615 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				14683 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				14719 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				14764 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				14812 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				14855 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				14860 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				14885 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				14888 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				14917 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				14919 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				14954 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				14956 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				15000 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				15023 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				15030 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				15053 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				15091 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				15125 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				15233 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				15254 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				15318 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				15686 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				15734 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				15817 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				15847 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				15855 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				15951 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				15975 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				15977 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				16000 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				16003 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				16021 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				16041 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				16154 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				16170 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				16174 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				16199 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				16215 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				16361 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				16386 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				16412 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				16439 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				16485 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				16543 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				16568 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				16572 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				16682 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				16687 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				16713 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				16717 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				16887 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				16925 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				17000 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				17017 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				17048 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				17053 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				17106 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				17192 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				17311 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				17320 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				17346 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				17359 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				17456 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				17498 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				17506 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				17584 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				17594 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				17607 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				17642 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				17643 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				17665 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				17681 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				17687 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				17696 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				17699 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				17705 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				17730 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				17732 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				17859 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				17861 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				18004 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				18011 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				18035 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				18054 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				18105 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				18107 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				18130 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				18173 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				18245 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				18269 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				18301 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				18327 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				18347 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				18620 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				18648 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				18660 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				18891 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				18934 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				18940 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				18959 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				18962 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				18969 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				18973 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				18977 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				19002 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				19085 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				19093 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				19150 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				19181 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				19257 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				19274 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				19289 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				19293 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				19385 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				19421 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				19455 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				19463 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				19477 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				19587 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				19625 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				19730 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				19754 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				19898 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				19933 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				20029 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				20086 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				20098 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				20117 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				20145 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				20161 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				20262 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				20287 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				20310 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				20322 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				20349 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				20384 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				20399 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				20461 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				20482 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				20523 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				20539 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				20550 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				20585 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				20677 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				20682 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				20711 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				20749 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				20874 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				20938 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				20941 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				21118 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				21119 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				21151 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				21183 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				21202 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				21265 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				21281 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				21300 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				21303 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				21312 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				21315 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				21416 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				21427 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				21487 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				21503 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				21531 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				21546 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				21631 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				21684 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				21705 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				21732 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				21755 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				21809 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				21862 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				21896 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				21924 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				21988 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				22001 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				22014 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				22057 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				22139 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				22143 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				22182 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				22204 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				22205 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				22258 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				22295 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				22346 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				22352 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				22397 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				22400 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				22409 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				22463 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				22562 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				22605 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				22647 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				22657 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				22666 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				22674 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				22677 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				22701 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				22706 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				22729 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				22785 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				22828 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				22833 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				22907 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				22915 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				22939 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				22950 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				22997 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				23021 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				23082 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				23099 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				23109 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				23129 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				23170 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				23209 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				23357 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				23371 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				23409 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				23431 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				23545 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				23557 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				23559 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				23573 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				23592 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				23666 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				23693 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				23721 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				23729 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				23844 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				23863 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				23870 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				23886 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				23986 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				23991 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				23994 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				24025 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				24042 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				24049 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				24096 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				24183 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				24196 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				24236 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				24275 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				24427 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				24461 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				24494 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				24501 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				24505 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				24506 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				24563 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				24568 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				24569 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				24616 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				24693 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				24694 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				24696 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				24703 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				24764 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				24799 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				24836 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				24849 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				24931 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				24943 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				24966 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				24985 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				24990 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				25079 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				25153 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				25156 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				25160 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				25185 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				25252 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				25311 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				25326 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				25474 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				25580 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				25584 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				25623 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				25678 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				25687 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				25768 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				25770 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				25917 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				25923 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				25943 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				25953 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				26031 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				26038 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				26083 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				26205 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				26332 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				26333 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				26335 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				26350 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				26352 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				26360 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				26366 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				26370 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				26411 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				26435 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				26537 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				26543 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				26628 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				26632 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				26642 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				26675 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				26795 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				26835 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				26844 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				26847 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				26855 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				26987 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				27078 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				27218 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				27249 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				27307 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				27366 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				27413 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				27500 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				27506 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				27585 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				27605 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				27658 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				27681 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				27725 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				27773 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				27831 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				27850 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				27862 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				27890 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				27902 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				27924 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				27930 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				27936 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				27955 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				28043 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				28105 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				28163 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				28229 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				28235 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				28247 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				28286 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				28331 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				28348 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				28371 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				28378 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				28433 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				28500 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				28517 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				28631 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				28695 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				28700 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				28713 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				28774 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				28791 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				28847 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				28850 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				28869 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				28889 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				28901 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				28904 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				28998 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				29082 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				29096 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				29120 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				29180 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				29238 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				29280 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				29371 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				29397 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				29478 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				29480 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				29504 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				29525 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				29621 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				29658 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				29670 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				29756 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				29770 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				29808 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				29818 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				29956 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				29964 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				29966 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				30025 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				30051 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				30081 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				30138 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				30164 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				30263 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				30317 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				30345 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				30354 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				30417 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				30482 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				30503 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				30702 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				30763 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				30789 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				30817 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				30823 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				30992 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				31041 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				31100 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				31111 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				31140 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				31172 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				31178 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				31300 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				31348 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				31424 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				31479 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				31503 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				31548 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				31564 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				31632 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				31645 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				31657 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				31671 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				31705 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				31736 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				31789 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				31801 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				31882 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				31896 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				31901 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				31903 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				31908 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				31960 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				31969 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				32017 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				32064 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				32091 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				32119 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				32126 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				32177 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				32250 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				32267 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				32392 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				32521 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				32572 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				32613 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				32684 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				32695 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				32754 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				32756 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				32766 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				32794 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				32832 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				32857 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				32939 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				32959 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				32987 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				33007 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				33018 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				33036 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				33058 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				33084 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				33090 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				33163 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				33166 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				33208 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				33277 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				33308 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				33311 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				33316 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				33367 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				33380 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				33494 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				33528 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				33580 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				33639 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				33646 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				33722 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				33726 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				33746 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				33787 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				33808 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				33843 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				33881 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				33917 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				34095 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				34146 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				34154 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				34186 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				34204 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				34216 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				34226 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				34290 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				34375 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				34379 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				34413 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				34458 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				34460 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				34502 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				34542 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				34559 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				34679 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				34683 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				34687 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				34709 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				34747 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				34749 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				34783 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				34802 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				34833 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				34850 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				34917 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				34999 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				35022 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				35056 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				35066 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				35091 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				35136 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				35211 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				35254 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				35255 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				35325 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				35378 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				35397 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				35472 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				35524 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				35562 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				35568 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				35580 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				35625 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				35682 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				35787 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				35819 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				35840 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				35869 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				35903 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				35904 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				36011 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				36030 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				36034 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				36039 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				36108 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				36172 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				36254 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				36261 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				36267 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				36285 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				36347 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				36377 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				36395 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				36490 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				36510 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				36626 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				36739 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				36758 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				36780 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				36839 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				36849 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				36888 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				36918 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				36926 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				36929 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				36994 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				37025 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				37053 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				37113 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				37159 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				37257 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				37287 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				37316 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				37330 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				37334 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				37336 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				37372 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				37446 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				37468 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				37479 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				37495 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				37499 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				37635 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				37717 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				37816 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				37929 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				37939 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				37961 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				38038 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				38039 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				38051 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				38091 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				38184 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				38189 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				38219 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				38220 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				38316 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				38344 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				38391 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				38466 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				38488 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				38502 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				38507 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				38591 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				38617 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				38620 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				38624 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				38637 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				38671 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				38676 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				38743 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				38773 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				38805 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				38834 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				38844 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				38902 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				38975 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				39030 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				39034 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				39043 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				39051 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				39055 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				39076 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				39090 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				39124 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				39147 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				39308 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				39327 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				39368 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				39372 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				39432 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				39455 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				39482 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				39525 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				39568 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				39569 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				39586 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				39598 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				39632 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				39673 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				39674 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				39676 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				39730 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				39755 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				39773 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				39805 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				39822 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				39828 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				39843 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				39849 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				39867 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				39951 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				39954 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				40029 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				40046 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				40094 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				40166 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				40185 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				40209 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				40222 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				40236 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				40270 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				40271 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				40277 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				40288 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				40302 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				40343 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				40359 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				40365 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				40385 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				40420 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				40430 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				40431 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				40451 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				40463 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				40476 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				40489 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				40492 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				40524 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				40530 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				40547 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				40568 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				40572 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				40601 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				40791 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				40798 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				40820 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				40863 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				40866 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				40867 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				40878 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				40895 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				40941 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				40966 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				40983 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				41010 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				41025 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				41047 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				41048 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				41143 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				41187 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				41215 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				41243 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				41335 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				41379 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				41429 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				41465 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				41527 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				41558 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				41569 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				41571 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				41600 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				41631 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				41857 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				41865 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				41909 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				41916 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				41940 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				41984 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				42118 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				42203 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				42221 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				42224 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				42227 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				42248 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				42351 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				42366 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				42367 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				42371 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				42504 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				42562 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				42686 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				42689 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				42717 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				42747 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				42774 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				42793 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				42808 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				42844 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				42855 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				42896 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				42909 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				42950 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				42981 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				43019 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				43083 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				43178 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				43197 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				43350 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				43354 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				43364 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				43375 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				43406 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				43436 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				43516 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				43588 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				43626 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				43648 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				43649 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				43725 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				43781 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				43809 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				43867 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				43908 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				43921 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				43934 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				43990 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				43995 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				44071 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				44216 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				44271 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				44364 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				44387 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				44432 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				44459 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				44470 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				44503 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				44533 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				44586 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				44656 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				44670 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				44676 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				44698 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				44706 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				44712 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				44734 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				44768 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				44793 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				44797 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				44823 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				44833 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				44838 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				44842 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				44851 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				44900 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				44915 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				44919 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				44938 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				44953 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				44958 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				44971 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				44998 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				45116 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				45174 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				45195 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				45256 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				45285 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				45441 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				45447 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				45472 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				45646 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				45656 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				45662 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				45820 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				45862 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				45887 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				45982 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				46014 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				46023 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				46075 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				46112 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				46138 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				46139 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				46207 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				46211 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				46230 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				46304 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				46372 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				46394 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				46437 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				46493 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				46496 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				46580 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				46636 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				46708 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				46733 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				46772 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				46783 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				46800 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				46828 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				46946 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				46986 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				46990 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				46999 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				47030 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				47109 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				47146 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				47172 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				47184 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				47194 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				47215 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				47239 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				47277 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				47442 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				47532 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				47597 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				47608 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				47715 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				47724 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				47727 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				47742 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				47748 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				47775 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				47801 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				47839 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				47937 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				47946 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				47980 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				48011 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				48065 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				48087 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				48103 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				48217 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				48253 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				48256 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				48291 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				48301 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				48325 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				48416 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				48565 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				48665 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				48675 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				48754 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				48793 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				48806 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				48849 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				48864 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				48888 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				48896 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				48905 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				49053 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				49081 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				49088 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				49089 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				49152 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				49225 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				49246 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				49251 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				49283 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				49293 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				49299 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				49390 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				49417 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				49510 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				49513 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				49531 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				49713 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				49737 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				49768 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				49772 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				49787 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				49812 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				49839 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				49841 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				49847 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				49870 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				49871 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				49902 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				49903 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				49956 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				49992 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				50183 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				50262 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				50356 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				50363 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				50443 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				50449 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				50481 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				50522 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				50543 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				50554 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				50570 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				50584 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				50627 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				50664 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				50849 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				50928 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				51006 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				51011 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				51040 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				51078 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				51106 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				51259 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				51308 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				51351 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				51352 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				51496 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				51502 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				51629 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				51682 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				51731 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				51778 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				51816 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				51820 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				51839 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				51950 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				52027 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				52039 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				52072 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				52304 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				52312 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				52368 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				52411 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				52468 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				52498 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				52530 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				52613 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				52631 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				52657 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				52665 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				52695 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				52714 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				52756 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				52786 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				52788 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				52908 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				52956 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				52981 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				53012 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				53088 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				53089 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				53265 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				53267 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				53302 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				53304 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				53309 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				53321 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				53329 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				53411 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				53499 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				53503 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				53536 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				53546 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				53568 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				53616 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				53622 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				53638 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				53658 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				53676 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				53791 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				53793 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				53794 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				53824 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				53852 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				53971 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				53996 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				54082 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				54124 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				54167 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				54170 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				54172 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				54221 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				54297 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				54298 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				54323 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				54340 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				54415 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				54557 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				54579 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				54594 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				54596 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				54606 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				54703 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				54715 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				54748 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				54813 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				54862 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				54929 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				54950 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				54957 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				55011 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				55041 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				55078 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				55160 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				55235 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				55256 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				55308 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				55317 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				55371 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				55394 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				55506 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				55510 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				55548 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				55560 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				55622 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				55761 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				55768 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				55825 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				55848 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				55864 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				55888 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				55893 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				55899 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				56029 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				56047 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				56100 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				56135 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				56142 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				56161 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				56188 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				56264 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				56340 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				56410 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				56445 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				56498 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				56519 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				56557 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				56589 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				56650 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				56651 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				56701 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				56712 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				56765 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				56783 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				56975 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				56993 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				57014 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				57031 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				57047 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				57074 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				57215 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				57233 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				57240 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				57246 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				57250 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				57346 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				57406 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				57412 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				57451 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				57492 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				57505 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				57509 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				57515 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				57609 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				57680 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				57683 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				57710 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				57716 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				57777 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				57867 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				57884 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				57974 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				58014 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				58017 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				58027 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				58032 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				58033 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				58119 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				58126 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				58230 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				58412 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				58449 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				58513 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				58519 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				58602 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				58630 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				58657 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				58679 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				58695 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				58830 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				58868 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				58939 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				58949 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				58961 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				58979 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				58997 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				59062 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				59077 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				59102 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				59117 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				59173 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				59211 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				59227 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				59262 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				59268 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				59275 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				59298 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				59310 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				59328 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				59347 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				59420 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				59491 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				59506 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				59556 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				59558 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				59574 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				59675 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				59720 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				59770 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				59772 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				59800 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				59871 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				59879 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				59881 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				59885 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				59887 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				59948 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				60000 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				60001 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				60065 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				60090 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				60102 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				60232 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				60297 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				60323 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				60328 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				60425 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				60426 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				60437 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				60460 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				60536 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				60578 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				60632 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				60664 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				60708 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				60765 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				60774 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				60793 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				60884 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				60930 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				60947 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				60951 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				60966 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				61036 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				61042 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				61090 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				61096 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				61101 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				61135 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				61169 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				61279 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				61310 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				61414 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				61464 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				61468 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				61482 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				61501 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				61511 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				61514 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				61516 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				61536 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				61544 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				61560 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				61577 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				61593 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				61644 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				61657 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				61680 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				61718 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				61742 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				61749 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				61773 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				61840 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				61874 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				61972 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				62009 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				62052 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				62062 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				62136 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				62144 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				62163 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				62192 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				62194 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				62275 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				62280 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				62300 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				62346 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				62379 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				62383 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				62449 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				62546 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				62548 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				62598 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				62603 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				62624 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				62750 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				62765 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				62785 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				62820 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				62835 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				62840 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				62846 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				62850 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				62893 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				62895 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				62943 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				62989 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				63013 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				63046 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				63092 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				63134 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				63142 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				63218 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				63233 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				63235 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				63279 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				63303 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				63305 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				63327 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				63332 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				63363 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				63409 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				63474 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				63477 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				63566 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				63571 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				63586 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				63615 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				63619 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				63663 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				63732 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				63767 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				63769 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				63868 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				63921 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				63947 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				63986 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				64010 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				64024 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				64029 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				64062 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				64095 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				64099 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				64120 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				64196 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				64294 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				64299 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				64328 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				64342 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				64345 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				64404 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				64455 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				64472 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				64475 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				64487 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				64497 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				64545 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				64560 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				64573 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				64649 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				64684 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				64696 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				64779 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				64855 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				64863 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				64900 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				64967 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				64990 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				65005 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				65017 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				65073 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				65102 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				65293 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				65344 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				65378 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				65382 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				65397 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				65399 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				65434 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				65491 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				65533 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),

                                OTHERS => STD_LOGIC_VECTOR(to_unsigned(99, 8))
                            );
                    
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
                ASSERT (mem_we = '1' OR mem_we = '0') REPORT "o_mem_we in an unexpected state" SEVERITY failure;
            END IF;
            ASSERT (enable_wire = '1' OR enable_wire = '0') REPORT "o_mem_en in an unexpected state" SEVERITY failure;
        END IF;
    END PROCESS;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    createScenario : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '0' THEN
            tb_rst <= scenario_rst(0);
            tb_w <= scenario_w(0);
            tb_start <= scenario_start(0);
            scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_done = '0' REPORT "TEST FALLITO (postreset DONE != 0 )" SEVERITY failure;
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(99, 8)) severity failure; --0001100111011101:99
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(99, 8)) severity failure; --1001010011101101:99
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z2 = std_logic_vector(to_unsigned(99, 8)) severity failure; --10101011001:99
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(99, 8)) severity failure; --010101111010001:99
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(99, 8)) severity failure; --1101000101001001:99
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(99, 8)) severity failure; --10100101111011:99
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(99, 8)) severity failure; --11101111001:99
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(99, 8)) severity failure; --10100101100101:99
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(99, 8)) severity failure; --10110001111011:99
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z1 = std_logic_vector(to_unsigned(99, 8)) severity failure; --000110011100011:99
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 

        ASSERT false REPORT "Simulation Ended! TEST PASSATO (EXAMPLE)" SEVERITY failure;
    END PROCESS testRoutine;

END projecttb;
