LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 1237; 
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00110" & "00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000" & "11111111111111111000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000011111111111111111000000000000000111111111111111100000000000011111111111111111100000000000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000001111111111111111100000000000000111111111111111111000000011111111111111111100000000011111111111111110000000000000000000000000000000111111111111111111000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000000011111111111111111000000000000000000000000000000111111111111111111000000000000011111111111111110000000000000000000011111111111111111100000000000000000000000000000001111111111111111110000000000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000000000001111111111111111110000000000000000000000000000000111111111111111111000000000011111111111110000000000111111111111111111000000000000000000000000000000011111111111111111100000000000000000000000000000011111111111111111100000000000000000000000000011111111111111000000000000000111111111111111110000000000000000000000000";
    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000" & "11110001111010001000000000000000000000010010101001100100000000000000000000000010000001100100000000000000000000000001110011010110110100000000000000000000000000010110001111100110000000000000000111001001101010100000000000001111110100101000100000000000000000000000000010111011110100011000000000000000000000001110011010001101000000000000000000111000111000010100000000000000011100110001000100000000000111000100100010000000000000111100111010000000000000000000000000000000000101011001111011110000000000000100010000111000000000000000000000000001010011110110000100000000000000000000001011111010001010010000000000000000000000000000001110100011001111000000000000000000000000000000001001010011111001000000000000011110000111010000000000000000000000011101011000001111100000000000000000000000000000000011011101000100000000000000000000000000000000001111010100000100100000000000000000000000110011000001111000000000000000000000000000000001110100011110110110000000000000000000000000000000111011000000101011000000000001110010010110000000000111111111100001001000000000000000000000000000000011100011000100001100000000000000000000000000000010111110110101100100000000000000000000000000011100101110101000000000000000011010010011011010000000000000000000000000";

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (  
				2 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				7 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				49 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				60 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				84 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				113 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				190 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				256 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				322 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				330 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				348 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				365 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				402 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				424 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				426 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				437 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				454 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				485 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				492 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				516 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				557 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				595 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				607 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				698 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				724 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				747 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				752 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				846 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				875 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				908 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				914 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				952 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				967 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				978 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				999 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				1082 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				1096 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				1122 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				1127 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				1163 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				1246 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				1258 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				1300 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				1317 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				1335 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				1345 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				1371 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				1392 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				1505 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				1559 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				1613 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				1647 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				1808 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				1857 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				1956 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				2046 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				2058 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				2060 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				2081 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				2160 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				2176 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				2304 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				2338 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				2358 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				2359 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				2425 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				2426 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				2441 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				2497 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				2504 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				2527 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				2573 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				2607 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				2616 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				2621 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				2697 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				2804 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				2850 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				2955 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				2956 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				2981 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				3080 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				3129 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				3137 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				3161 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				3170 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				3231 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				3253 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				3261 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				3267 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				3308 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				3320 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				3329 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				3379 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				3397 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				3493 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				3535 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				3611 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				3627 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				3633 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				3673 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				3675 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				3686 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				3699 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				3738 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				3742 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				3758 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				3822 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				3851 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				3883 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				4062 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				4083 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				4091 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				4098 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				4100 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				4142 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				4342 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				4349 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				4400 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				4423 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				4439 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				4460 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				4463 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				4474 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				4479 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				4480 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				4498 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				4626 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				4640 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				4662 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				4681 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				4683 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				4720 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				4744 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				4755 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				4766 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				4806 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				4832 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				4861 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				4876 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				4957 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				4964 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				5134 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				5174 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				5200 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				5206 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				5208 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				5221 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				5224 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				5257 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				5297 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				5325 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				5330 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				5333 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				5357 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				5362 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				5383 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				5399 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				5467 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				5479 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				5593 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				5661 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				5666 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				5669 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				5745 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				5780 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				5836 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				5852 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				5907 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				5910 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				5922 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				5926 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				5945 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				5983 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				5988 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				6064 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				6142 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				6185 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				6276 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				6339 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				6352 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				6382 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				6403 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				6468 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				6497 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				6528 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				6573 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				6578 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				6607 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				6667 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				6684 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				6731 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				6954 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				6955 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				6966 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				6974 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				6987 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				7063 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				7093 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				7121 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				7122 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				7185 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				7203 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				7214 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				7247 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				7310 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				7352 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				7353 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				7358 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				7359 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				7431 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				7459 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				7472 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				7508 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				7526 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				7533 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				7536 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				7539 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				7609 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				7640 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				7655 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				7681 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				7733 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				7813 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				7873 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				7915 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				8148 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				8181 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				8187 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				8272 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				8332 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				8365 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				8476 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				8538 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				8602 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				8621 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				8659 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				8670 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				8768 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				8793 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				8800 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				8830 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				8941 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				8978 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				8999 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				9027 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				9178 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				9188 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				9239 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				9266 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				9283 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				9296 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				9342 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				9453 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				9459 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				9509 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				9536 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				9541 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				9573 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				9577 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				9594 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				9604 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				9658 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				9695 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				9734 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				9747 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				9807 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				9838 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				9843 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				9894 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				9936 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				9969 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				9970 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				9990 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				10018 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				10047 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				10055 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				10057 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				10107 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				10126 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				10132 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				10205 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				10239 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				10347 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				10359 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				10414 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				10445 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				10537 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				10607 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				10691 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				10698 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				10741 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				10744 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				10754 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				10782 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				10784 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				10808 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				10813 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				10923 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				10926 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				10933 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				10946 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				11114 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				11127 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				11212 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				11234 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				11238 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				11239 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				11279 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				11327 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				11339 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				11474 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				11609 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				11710 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				11730 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				11737 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				11742 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				11772 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				11797 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				11822 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				11836 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				11837 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				11840 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				11861 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				11864 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				11906 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				12020 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				12027 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				12066 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				12100 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				12120 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				12178 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				12195 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				12209 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				12248 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				12260 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				12303 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				12315 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				12344 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				12365 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				12370 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				12372 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				12376 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				12495 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				12533 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				12618 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				12658 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				12667 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				12704 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				12734 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				12741 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				12755 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				12794 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				12920 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				12968 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				12976 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				13005 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				13014 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				13048 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				13097 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				13125 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				13153 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				13159 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				13161 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				13221 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				13316 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				13326 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				13411 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				13431 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				13473 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				13485 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				13537 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				13616 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				13637 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				13680 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				13703 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				13782 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				13807 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				13876 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				13879 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				13882 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				13897 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				13947 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				13969 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				13978 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				14028 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				14055 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				14109 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				14207 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				14212 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				14266 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				14284 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				14288 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				14360 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				14367 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				14425 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				14430 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				14473 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				14508 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				14515 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				14587 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				14622 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				14700 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				14731 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				14738 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				14741 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				14745 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				14812 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				14848 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				14897 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				14899 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				14942 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				14960 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				15008 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				15082 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				15110 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				15115 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				15121 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				15183 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				15281 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				15305 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				15358 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				15373 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				15427 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				15462 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				15514 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				15515 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				15584 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				15677 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				15686 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				15708 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				15738 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				15789 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				15823 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				15884 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				15933 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				15975 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				16005 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				16110 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				16152 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				16247 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				16305 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				16312 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				16349 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				16380 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				16383 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				16412 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				16429 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				16483 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				16484 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				16514 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				16583 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				16586 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				16647 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				16659 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				16763 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				16783 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				16788 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				16967 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				17137 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				17211 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				17256 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				17258 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				17276 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				17278 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				17284 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				17297 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				17308 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				17342 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				17360 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				17369 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				17398 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				17412 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				17500 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				17514 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				17542 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				17749 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				17764 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				17796 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				17809 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				17837 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				17919 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				17975 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				18053 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				18235 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				18251 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				18304 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				18305 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				18352 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				18370 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				18422 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				18459 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				18566 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				18600 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				18619 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				18652 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				18700 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				18712 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				18768 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				18785 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				18802 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				18843 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				18949 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				18997 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				19095 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				19127 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				19137 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				19144 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				19159 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				19170 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				19172 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				19180 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				19212 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				19245 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				19271 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				19280 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				19301 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				19309 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				19367 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				19398 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				19546 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				19561 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				19579 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				19580 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				19639 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				19660 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				19667 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				19725 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				19730 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				19765 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				19784 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				19848 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				19849 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				19872 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				19874 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				19881 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				19933 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				19951 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				19978 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				20045 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				20078 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				20157 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				20158 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				20191 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				20282 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				20357 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				20394 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				20417 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				20433 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				20438 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				20525 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				20526 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				20640 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				20661 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				20684 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				20738 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				20767 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				20807 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				20850 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				20953 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				21016 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				21029 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				21077 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				21131 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				21154 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				21182 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				21255 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				21341 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				21583 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				21587 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				21600 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				21769 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				21796 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				21813 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				21905 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				21996 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				22035 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				22066 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				22124 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				22142 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				22239 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				22279 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				22349 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				22385 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				22402 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				22484 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				22486 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				22537 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				22567 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				22579 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				22593 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				22624 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				22652 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				22656 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				22657 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				22712 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				22745 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				22752 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				22834 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				22924 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				22956 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				23020 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				23032 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				23041 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				23054 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				23096 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				23105 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				23153 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				23205 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				23214 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				23290 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				23373 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				23442 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				23444 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				23455 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				23461 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				23481 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				23485 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				23525 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				23601 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				23618 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				23619 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				23661 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				23843 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				23876 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				23878 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				23889 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				23973 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				24025 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				24091 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				24100 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				24103 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				24128 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				24170 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				24185 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				24199 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				24220 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				24223 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				24229 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				24232 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				24269 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				24366 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				24383 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				24398 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				24451 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				24456 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				24519 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				24537 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				24542 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				24546 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				24583 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				24609 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				24614 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				24618 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				24729 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				24839 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				24845 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				24912 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				25018 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				25025 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				25035 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				25066 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				25127 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				25166 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				25268 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				25298 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				25338 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				25565 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				25616 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				25644 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				25688 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				25763 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				25769 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				25862 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				25877 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				25883 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				25889 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				25891 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				25902 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				26008 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				26074 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				26160 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				26185 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				26196 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				26210 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				26281 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				26289 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				26328 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				26367 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				26376 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				26440 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				26446 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				26451 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				26494 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				26521 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				26547 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				26577 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				26586 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				26593 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				26614 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				26633 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				26687 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				26784 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				26822 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				26838 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				26871 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				26890 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				26931 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				26944 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				26962 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				26971 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				26991 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				27018 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				27068 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				27080 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				27092 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				27126 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				27189 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				27239 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				27257 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				27274 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				27280 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				27329 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				27342 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				27419 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				27426 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				27490 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				27508 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				27536 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				27549 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				27610 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				27630 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				27643 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				27661 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				27667 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				27740 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				27795 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				27797 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				27806 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				27840 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				27873 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				28022 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				28061 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				28134 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				28272 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				28296 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				28311 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				28326 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				28329 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				28333 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				28456 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				28477 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				28490 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				28511 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				28525 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				28538 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				28574 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				28591 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				28617 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				28733 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				28743 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				28788 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				28881 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				28886 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				28915 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				28939 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				28953 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				28960 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				28970 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				29030 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				29047 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				29113 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				29120 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				29133 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				29136 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				29228 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				29263 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				29265 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				29315 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				29334 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				29393 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				29394 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				29481 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				29491 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				29509 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				29519 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				29523 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				29527 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				29543 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				29570 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				29589 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				29612 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				29655 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				29665 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				29691 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				29694 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				29704 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				29780 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				29800 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				29900 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				29918 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				29921 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				29928 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				30018 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				30020 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				30036 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				30049 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				30050 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				30123 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				30141 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				30196 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				30206 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				30214 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				30244 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				30268 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				30269 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				30331 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				30345 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				30387 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				30438 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				30468 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				30559 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				30561 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				30582 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				30629 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				30671 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				30676 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				30753 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				30762 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				30765 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				30826 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				30835 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				30843 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				30879 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				30898 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				30934 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				31035 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				31051 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				31106 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				31168 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				31180 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				31202 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				31214 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				31239 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				31289 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				31305 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				31332 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				31381 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				31383 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				31411 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				31476 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				31488 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				31519 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				31535 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				31585 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				31599 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				31615 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				31646 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				31673 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				31766 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				31775 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				31776 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				31796 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				31799 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				31801 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				31838 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				31857 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				31865 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				31964 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				32002 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				32021 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				32031 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				32036 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				32115 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				32203 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				32212 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				32437 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				32519 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				32529 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				32554 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				32626 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				32659 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				32676 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				32710 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				32722 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				32821 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				32852 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				32871 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				32918 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				32990 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				33023 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				33053 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				33099 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				33105 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				33157 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				33179 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				33185 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				33254 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				33299 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				33322 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				33355 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				33371 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				33373 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				33442 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				33453 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				33513 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				33610 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				33663 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				33714 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				33735 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				33854 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				33867 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				33957 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				33968 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				34014 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				34048 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				34066 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				34080 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				34103 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				34156 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				34178 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				34213 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				34214 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				34238 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				34331 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				34362 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				34374 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				34378 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				34386 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				34427 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				34473 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				34493 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				34515 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				34555 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				34657 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				34698 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				34709 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				34710 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				34718 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				34738 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				34825 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				34827 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				34868 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				34871 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				34873 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				34903 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				34905 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				34933 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				34999 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				35022 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				35038 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				35121 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				35151 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				35153 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				35215 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				35272 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				35273 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				35283 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				35285 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				35293 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				35297 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				35316 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				35324 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				35326 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				35328 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				35363 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				35492 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				35493 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				35500 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				35561 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				35654 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				35668 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				35728 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				35744 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				36066 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				36129 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				36209 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				36225 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				36400 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				36417 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				36448 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				36501 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				36506 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				36529 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				36536 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				36539 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				36558 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				36559 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				36611 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				36675 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				36702 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				36704 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				36761 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				36830 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				36832 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				36880 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				36916 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				36920 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				36933 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				36945 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				36962 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				36977 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				37017 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				37029 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				37045 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				37072 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				37121 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				37138 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				37259 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				37298 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				37332 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				37420 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				37482 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				37571 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				37598 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				37664 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				37687 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				37728 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				37830 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				37856 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				37870 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				37907 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				37960 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				37971 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				38009 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				38050 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				38109 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				38112 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				38189 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				38203 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				38230 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				38231 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				38280 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				38282 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				38306 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				38393 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				38414 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				38463 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				38524 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				38538 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				38543 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				38584 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				38663 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				38666 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				38746 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				38890 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				38902 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				38956 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				38958 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				38987 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				39001 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				39020 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				39026 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				39046 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				39188 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				39209 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				39310 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				39342 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				39346 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				39378 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				39494 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				39502 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				39517 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				39570 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				39573 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				39595 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				39602 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				39659 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				39753 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				39869 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				39881 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				39962 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				39964 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				39990 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				40009 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				40071 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				40108 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				40135 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				40145 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				40175 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				40237 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				40264 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				40324 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				40326 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				40388 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				40457 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				40551 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				40556 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				40561 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				40575 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				40624 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				40688 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				40711 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				40712 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				40723 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				40764 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				40794 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				40853 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				40975 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				41003 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				41025 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				41105 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				41134 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				41162 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				41201 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				41205 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				41231 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				41245 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				41263 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				41274 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				41280 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				41313 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				41338 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				41379 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				41421 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				41457 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				41471 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				41485 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				41511 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				41694 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				41726 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				41751 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				41820 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				41842 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				41883 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				41890 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				41899 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				42006 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				42011 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				42015 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				42017 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				42036 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				42053 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				42055 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				42139 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				42169 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				42202 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				42225 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				42226 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				42247 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				42338 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				42355 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				42478 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				42515 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				42560 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				42567 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				42584 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				42592 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				42690 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				42714 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				42715 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				42726 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				42748 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				42755 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				42781 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				42814 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				42825 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				42835 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				42837 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				42846 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				42859 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				42884 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				42950 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				42991 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				43057 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				43069 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				43205 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				43249 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				43252 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				43300 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				43368 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				43405 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				43430 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				43477 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				43481 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				43588 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				43634 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				43686 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				43711 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				43829 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				43869 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				43982 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				44019 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				44024 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				44032 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				44050 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				44171 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				44184 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				44251 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				44297 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				44317 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				44435 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				44448 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				44493 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				44494 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				44525 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				44578 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				44580 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				44609 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				44723 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				44735 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				44752 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				44883 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				44894 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				44913 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				44933 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				44945 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				45022 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				45098 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				45198 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				45210 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				45271 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				45281 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				45316 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				45318 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				45325 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				45389 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				45404 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				45411 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				45428 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				45432 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				45458 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				45463 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				45472 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				45563 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				45596 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				45613 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				45740 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				45868 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				45916 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				45956 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				45957 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				46001 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				46016 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				46037 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				46048 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				46159 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				46187 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				46218 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				46274 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				46275 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				46311 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				46327 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				46343 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				46347 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				46356 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				46384 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				46388 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				46392 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				46405 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				46421 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				46460 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				46568 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				46624 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				46649 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				46688 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				46706 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				46813 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				46845 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				47025 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				47120 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				47144 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				47151 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				47328 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				47348 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				47426 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				47432 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				47486 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				47632 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				47647 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				47692 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				47720 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				47735 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				47759 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				47779 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				47802 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				47805 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				47826 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				47872 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				47923 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				47947 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				47977 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				48088 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				48132 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				48163 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				48171 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				48224 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				48231 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				48233 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				48258 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				48265 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				48290 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				48333 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				48347 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				48349 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				48351 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				48352 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				48381 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				48416 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				48436 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				48460 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				48558 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				48596 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				48644 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				48696 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				48775 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				48786 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				48793 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				48796 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				48883 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				48889 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				48945 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				48972 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				48978 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				48996 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				49050 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				49129 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				49201 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				49258 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				49308 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				49318 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				49433 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				49476 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				49494 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				49498 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				49512 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				49581 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				49642 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				49668 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				49672 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				49703 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				49761 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				49765 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				49790 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				49828 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				49941 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				49959 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				50007 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				50035 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				50066 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				50090 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				50195 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				50199 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				50219 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				50239 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				50248 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				50279 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				50280 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				50281 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				50389 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				50432 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				50440 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				50491 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				50497 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				50568 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				50574 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				50649 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				50655 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				50692 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				50719 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				50729 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				50817 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				50831 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				50906 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				50918 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				50928 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				51025 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				51072 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				51087 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				51157 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				51158 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				51232 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				51259 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				51297 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				51407 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				51428 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				51446 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				51506 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				51516 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				51525 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				51527 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				51602 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				51621 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				51641 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				51670 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				51894 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				51922 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				52016 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				52102 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				52116 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				52141 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				52174 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				52184 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				52213 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				52225 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				52253 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				52288 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				52392 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				52461 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				52467 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				52486 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				52576 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				52625 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				52650 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				52673 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				52683 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				52696 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				52755 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				52759 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				52806 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				52834 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				52863 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				52870 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				52879 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				52984 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				53000 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				53014 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				53035 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				53058 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				53085 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				53158 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				53169 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				53189 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				53192 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				53250 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				53270 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				53299 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				53308 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				53341 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				53442 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				53468 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				53476 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				53505 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				53514 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				53590 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				53599 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				53604 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				53609 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				53627 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				53738 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				54059 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				54060 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				54062 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				54073 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				54200 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				54209 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				54226 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				54234 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				54278 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				54336 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				54352 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				54431 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				54433 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				54470 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				54603 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				54689 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				54710 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				54742 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				54785 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				54814 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				54910 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				54953 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				54957 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				54971 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				54987 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				55012 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				55151 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				55159 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				55166 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				55173 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				55262 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				55308 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				55312 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				55343 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				55347 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				55415 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				55565 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				55590 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				55666 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				55747 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				55878 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				55882 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				55883 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				55893 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				55936 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				55937 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				55992 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				56022 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				56024 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				56079 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				56085 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				56138 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				56144 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				56170 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				56235 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				56260 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				56289 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				56294 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				56364 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				56382 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				56394 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				56436 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				56437 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				56451 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				56475 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				56500 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				56612 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				56647 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				56759 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				56761 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				56770 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				56782 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				56808 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				56828 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				56882 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				56954 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				57026 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				57046 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				57085 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				57104 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				57109 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				57125 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				57168 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				57206 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				57217 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				57227 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				57258 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				57552 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				57559 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				57578 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				57586 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				57616 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				57665 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				57727 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				57739 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				57900 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				57910 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				58070 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				58073 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				58080 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				58084 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				58128 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				58198 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				58287 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				58331 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				58334 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				58366 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				58390 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				58394 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				58424 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				58461 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				58541 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				58558 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				58580 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				58630 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				58648 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				58654 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				58674 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				58770 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				58819 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				58863 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				58882 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				58897 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				58919 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				59035 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				59048 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				59182 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				59209 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				59240 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				59271 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				59321 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				59349 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				59370 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				59381 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				59436 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				59655 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				59702 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				59770 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				59827 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				59830 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				59864 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				59885 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				60023 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				60037 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				60048 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				60094 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				60123 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				60461 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				60468 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				60502 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				60515 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				60517 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				60553 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				60576 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				60601 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				60640 => STD_LOGIC_VECTOR(to_unsigned(255, 8)),
				60649 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				60680 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				60800 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				60823 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				60936 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				60951 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				61107 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				61138 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				61141 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				61165 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				61178 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				61196 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				61201 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				61232 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				61281 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				61316 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				61405 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				61415 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				61424 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				61439 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				61463 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				61489 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				61501 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				61539 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				61548 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				61555 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				61566 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				61604 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				61627 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				61640 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				61655 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				61709 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				61773 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				61935 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				61941 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				61951 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				61965 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				61999 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				62020 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				62044 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				62153 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				62173 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				62221 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				62224 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				62238 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				62282 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				62290 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				62293 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				62311 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				62448 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				62567 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				62584 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				62604 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				62613 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				62621 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				62636 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				62672 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				62694 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				62730 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				62737 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				62770 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				62835 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				62874 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				62896 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				62900 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				62925 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				62982 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				62999 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				63013 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				63040 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				63064 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				63073 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				63215 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				63238 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				63256 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				63291 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				63301 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				63311 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				63316 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				63318 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				63344 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				63364 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				63406 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				63445 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				63484 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				63503 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				63515 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				63517 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				63548 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				63686 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				63728 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				63753 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				63822 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				63877 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				63936 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				63965 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				64048 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				64079 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				64088 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				64096 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				64139 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				64151 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				64197 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				64200 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				64217 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				64245 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				64258 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				64259 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				64316 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				64327 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				64341 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				64369 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				64391 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				64437 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				64499 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				64500 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				64527 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				64538 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				64641 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				64668 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				64736 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				64775 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				64791 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				64811 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				64865 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				64876 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				64890 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				64977 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				64982 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				65053 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				65095 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				65112 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				65137 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				65259 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				65279 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				65353 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				65426 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				65432 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				65457 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				65493 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				65497 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),

                                OTHERS => STD_LOGIC_VECTOR(to_unsigned(231, 8))
                            );
                    
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
                ASSERT (mem_we = '1' OR mem_we = '0') REPORT "o_mem_we in an unexpected state" SEVERITY failure;
            END IF;
            ASSERT (enable_wire = '1' OR enable_wire = '0') REPORT "o_mem_en in an unexpected state" SEVERITY failure;
        END IF;
    END PROCESS;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    createScenario : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '0' THEN
            tb_rst <= scenario_rst(0);
            tb_w <= scenario_w(0);
            tb_start <= scenario_start(0);
            scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_done = '0' REPORT "TEST FALLITO (postreset DONE != 0 )" SEVERITY failure;
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 110001111010001:231->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1001010100110010:231->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 100000011001000:231->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1001101011011010:231->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 110001111100110:231->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 10010011010101:231->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1111101001010001:231->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 111011110100011:231->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 10011010001101:231->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 110001110000101:231->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1100110001000100:231->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1110001001000100:231->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 11110011101000:231->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1011001111011110:231->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1000100001110000:231->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1001111011000010:231->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1111101000101001:231->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 110100011001111:231->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1001010011111001:231->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 11000011101000:231->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1010110000011111:231->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1101110100010000:231->0 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 110101000001001:231->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 100110000011110:231->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1010001111011011:231->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1011000000101011:231->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 11001001011:231->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1111111100001001:231->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1000110001000011:231->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 1111101101011001:231->2 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 100101110101:231->3 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_start = '1';

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
	WAIT UNTIL tb_done = '1';
	WAIT FOR CLOCK_PERIOD/2;
	ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- 101001001101101:231->1 
	ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8)) severity failure; -- NOT UPDATED 
	WAIT UNTIL tb_done = '0';
	WAIT FOR CLOCK_PERIOD/2;

	ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
	ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
	ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
	ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 

        ASSERT false REPORT "Simulation Ended! TEST PASSATO (EXAMPLE)" SEVERITY failure;
    END PROCESS testRoutine;

END projecttb;